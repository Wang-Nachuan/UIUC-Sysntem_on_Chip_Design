
-------------------------------------------------------------------------------
-- VHDL test file for 'image.vhd'
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;
use std.env.stop;

entity image_test is
    generic(TREE_RAM_BITS: positive := 13;
            NUM_CLASSES:   positive := 2;
            NUM_FEATURES:  positive := 8);
end image_test;

architecture behavior of image_test is

    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;

             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);

             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;

             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;

    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;

    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto 0);
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';

    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);

    -- Clock period definition
    constant Clk_period : time := 10 ns;

    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');

    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

    -------------------- Newly added signals --------------------

    -- signal addr_count, addr_count_n: std_logic_vector(TREE_RAM_BITS - 1 downto 0);
    shared variable v_TIME : time := 0 ns;

begin

    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);

    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);

    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);

    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;

    -- Stimulus process
    stim_proc: process
    begin

        Reset <= '1';
        Addr <= "0000000000000";

        -- hold reset state for 100 ns.
        wait for 100 ns;

        Reset <= '0';

        wait for Clk_period*10;


-- LOAD TREES START
-----------------------------------------------------------------------

-- Class number = 2
-- Max depth = 7
-- Min depth = 7
-- Tree number = 12
-- average stand deviation for each class is: 
-- class 0 = 0.0
-- class 1 = 0.0

-- LOAD TREES
-----------------------------------------------------------------------

-- Load and valid trees flags
Load_trees <= '1';
Valid_node <= '1';

-- load tree numbers 
Addr <= "0000000000000";
Trees_din <= x"0000000c";
wait for Clk_period;

-- Reset load flag
Load_trees <= '0';    
    
-- Load starting address
--tree 0 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000001";
Trees_din <= "00000000000000000000000000001101";
wait for Clk_period;

--tree 1 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000010";
Trees_din <= "00000000000000000000000010001100";
wait for Clk_period;

--tree 2 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000011";
Trees_din <= "00000000000000000000000100001011";
wait for Clk_period;

--tree 3 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000100";
Trees_din <= "00000000000000000000000110001010";
wait for Clk_period;

--tree 4 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000101";
Trees_din <= "00000000000000000000001000001001";
wait for Clk_period;

--tree 5 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000110";
Trees_din <= "00000000000000000000001010001000";
wait for Clk_period;

--tree 6 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000000111";
Trees_din <= "00000000000000000010001100000111";
wait for Clk_period;

--tree 7 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000001000";
Trees_din <= "00000000000000000010001110000110";
wait for Clk_period;

--tree 8 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000001001";
Trees_din <= "00000000000000000010010000000101";
wait for Clk_period;

--tree 9 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000001010";
Trees_din <= "00000000000000000010010010000100";
wait for Clk_period;

--tree 10 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000001011";
Trees_din <= "00000000000000000010010100000011";
wait for Clk_period;

--tree 11 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000001100";
Trees_din <= "00000000000000000010010110000010";
wait for Clk_period;




----------tree 0-------------------

Addr <= "0000000001101";
Trees_din <= "00000010000000000000010110000000";
wait for Clk_period;
Addr <= "0000000001110";
Trees_din <= "00000011000000000100101101000000";
wait for Clk_period;
Addr <= "0000000001111";
Trees_din <= "00000010000000000001000000100000";
wait for Clk_period;
Addr <= "0000000010000";
Trees_din <= "00000000000000000011101100010000";
wait for Clk_period;
Addr <= "0000000010001";
Trees_din <= "00000011000000000110001100001000";
wait for Clk_period;
Addr <= "0000000010010";
Trees_din <= "00000111000000000001001100000100";
wait for Clk_period;
Addr <= "0000000010011";
Trees_din <= "00000000000100110000001000110001";
wait for Clk_period;
Addr <= "0000000010100";
Trees_din <= "00000000000111000000001000110001";
wait for Clk_period;
Addr <= "0000000010101";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0000000010110";
Trees_din <= "00000000010001110000001000110001";
wait for Clk_period;
Addr <= "0000000010111";
Trees_din <= "00000000000000100000001000110001";
wait for Clk_period;
Addr <= "0000000011000";
Trees_din <= "00000010000000000100101000001000";
wait for Clk_period;
Addr <= "0000000011001";
Trees_din <= "00000101000000000011100000000100";
wait for Clk_period;
Addr <= "0000000011010";
Trees_din <= "00000000010000000000001000110001";
wait for Clk_period;
Addr <= "0000000011011";
Trees_din <= "00000000011000100000001000110001";
wait for Clk_period;
Addr <= "0000000011100";
Trees_din <= "00000011000000000010100100000100";
wait for Clk_period;
Addr <= "0000000011101";
Trees_din <= "00000000001110100000001000110001";
wait for Clk_period;
Addr <= "0000000011110";
Trees_din <= "00000000001000100000001000110001";
wait for Clk_period;
Addr <= "0000000011111";
Trees_din <= "00000010000000000010110100010000";
wait for Clk_period;
Addr <= "0000000100000";
Trees_din <= "00000010000000000001000000001000";
wait for Clk_period;
Addr <= "0000000100001";
Trees_din <= "00000100000000000001010000000100";
wait for Clk_period;
Addr <= "0000000100010";
Trees_din <= "00000000010100100000001000110001";
wait for Clk_period;
Addr <= "0000000100011";
Trees_din <= "00000000010010000000001000110001";
wait for Clk_period;
Addr <= "0000000100100";
Trees_din <= "00000010000000000010111000000100";
wait for Clk_period;
Addr <= "0000000100101";
Trees_din <= "00000000001100000000001000110001";
wait for Clk_period;
Addr <= "0000000100110";
Trees_din <= "00000000001110110000001000110001";
wait for Clk_period;
Addr <= "0000000100111";
Trees_din <= "00000111000000000011111100001000";
wait for Clk_period;
Addr <= "0000000101000";
Trees_din <= "00000011000000000000101100000100";
wait for Clk_period;
Addr <= "0000000101001";
Trees_din <= "00000000000000010000001000110001";
wait for Clk_period;
Addr <= "0000000101010";
Trees_din <= "00000000000110000000001000110001";
wait for Clk_period;
Addr <= "0000000101011";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "0000000101100";
Trees_din <= "00000000001010010000001000110001";
wait for Clk_period;
Addr <= "0000000101101";
Trees_din <= "00000000000111100000001000110001";
wait for Clk_period;
Addr <= "0000000101110";
Trees_din <= "00000101000000000100010000100000";
wait for Clk_period;
Addr <= "0000000101111";
Trees_din <= "00000001000000000001100000010000";
wait for Clk_period;
Addr <= "0000000110000";
Trees_din <= "00000000000000000010011000001000";
wait for Clk_period;
Addr <= "0000000110001";
Trees_din <= "00000001000000000011001100000100";
wait for Clk_period;
Addr <= "0000000110010";
Trees_din <= "00000000000001110000001000110001";
wait for Clk_period;
Addr <= "0000000110011";
Trees_din <= "00000000010001010000001000110001";
wait for Clk_period;
Addr <= "0000000110100";
Trees_din <= "00000000000000000101000000000100";
wait for Clk_period;
Addr <= "0000000110101";
Trees_din <= "00000000010011110000001000110001";
wait for Clk_period;
Addr <= "0000000110110";
Trees_din <= "00000000000110000000001000110001";
wait for Clk_period;
Addr <= "0000000110111";
Trees_din <= "00000010000000000010011000001000";
wait for Clk_period;
Addr <= "0000000111000";
Trees_din <= "00000101000000000001000000000100";
wait for Clk_period;
Addr <= "0000000111001";
Trees_din <= "00000000001100110000001000110001";
wait for Clk_period;
Addr <= "0000000111010";
Trees_din <= "00000000001100100000001000110001";
wait for Clk_period;
Addr <= "0000000111011";
Trees_din <= "00000110000000000001100000000100";
wait for Clk_period;
Addr <= "0000000111100";
Trees_din <= "00000000000110010000001000110001";
wait for Clk_period;
Addr <= "0000000111101";
Trees_din <= "00000000001001000000001000110001";
wait for Clk_period;
Addr <= "0000000111110";
Trees_din <= "00000111000000000000001100010000";
wait for Clk_period;
Addr <= "0000000111111";
Trees_din <= "00000010000000000011101100001000";
wait for Clk_period;
Addr <= "0000001000000";
Trees_din <= "00000011000000000011100100000100";
wait for Clk_period;
Addr <= "0000001000001";
Trees_din <= "00000000000111010000001000110001";
wait for Clk_period;
Addr <= "0000001000010";
Trees_din <= "00000000010000110000001000110001";
wait for Clk_period;
Addr <= "0000001000011";
Trees_din <= "00000011000000000101011000000100";
wait for Clk_period;
Addr <= "0000001000100";
Trees_din <= "00000000011000110000001000110001";
wait for Clk_period;
Addr <= "0000001000101";
Trees_din <= "00000000000100110000001000110001";
wait for Clk_period;
Addr <= "0000001000110";
Trees_din <= "00000101000000000110000100001000";
wait for Clk_period;
Addr <= "0000001000111";
Trees_din <= "00000100000000000011111000000100";
wait for Clk_period;
Addr <= "0000001001000";
Trees_din <= "00000000010000010000001000110001";
wait for Clk_period;
Addr <= "0000001001001";
Trees_din <= "00000000001100110000001000110001";
wait for Clk_period;
Addr <= "0000001001010";
Trees_din <= "00000110000000000010110100000100";
wait for Clk_period;
Addr <= "0000001001011";
Trees_din <= "00000000001101000000001000110001";
wait for Clk_period;
Addr <= "0000001001100";
Trees_din <= "00000000001000110000001000110001";
wait for Clk_period;
Addr <= "0000001001101";
Trees_din <= "00000011000000000000111001000000";
wait for Clk_period;
Addr <= "0000001001110";
Trees_din <= "00000001000000000100101000100000";
wait for Clk_period;
Addr <= "0000001001111";
Trees_din <= "00000011000000000000000000010000";
wait for Clk_period;
Addr <= "0000001010000";
Trees_din <= "00000010000000000110000000001000";
wait for Clk_period;
Addr <= "0000001010001";
Trees_din <= "00000100000000000010011000000100";
wait for Clk_period;
Addr <= "0000001010010";
Trees_din <= "00000000000100010000001000110001";
wait for Clk_period;
Addr <= "0000001010011";
Trees_din <= "00000000010001000000001000110001";
wait for Clk_period;
Addr <= "0000001010100";
Trees_din <= "00000000000000000011001100000100";
wait for Clk_period;
Addr <= "0000001010101";
Trees_din <= "00000000010001010000001000110001";
wait for Clk_period;
Addr <= "0000001010110";
Trees_din <= "00000000001110000000001000110001";
wait for Clk_period;
Addr <= "0000001010111";
Trees_din <= "00000110000000000000001000001000";
wait for Clk_period;
Addr <= "0000001011000";
Trees_din <= "00000001000000000010101100000100";
wait for Clk_period;
Addr <= "0000001011001";
Trees_din <= "00000000000111010000001000110001";
wait for Clk_period;
Addr <= "0000001011010";
Trees_din <= "00000000000110010000001000110001";
wait for Clk_period;
Addr <= "0000001011011";
Trees_din <= "00000011000000000011101000000100";
wait for Clk_period;
Addr <= "0000001011100";
Trees_din <= "00000000010110100000001000110001";
wait for Clk_period;
Addr <= "0000001011101";
Trees_din <= "00000000001100100000001000110001";
wait for Clk_period;
Addr <= "0000001011110";
Trees_din <= "00000000000000000011100100010000";
wait for Clk_period;
Addr <= "0000001011111";
Trees_din <= "00000100000000000000010100001000";
wait for Clk_period;
Addr <= "0000001100000";
Trees_din <= "00000100000000000001010000000100";
wait for Clk_period;
Addr <= "0000001100001";
Trees_din <= "00000000000111110000001000110001";
wait for Clk_period;
Addr <= "0000001100010";
Trees_din <= "00000000001101110000001000110001";
wait for Clk_period;
Addr <= "0000001100011";
Trees_din <= "00000011000000000011001100000100";
wait for Clk_period;
Addr <= "0000001100100";
Trees_din <= "00000000000000000000001000110001";
wait for Clk_period;
Addr <= "0000001100101";
Trees_din <= "00000000010101010000001000110001";
wait for Clk_period;
Addr <= "0000001100110";
Trees_din <= "00000111000000000000101100001000";
wait for Clk_period;
Addr <= "0000001100111";
Trees_din <= "00000111000000000000111000000100";
wait for Clk_period;
Addr <= "0000001101000";
Trees_din <= "00000000010010010000001000110001";
wait for Clk_period;
Addr <= "0000001101001";
Trees_din <= "00000000010001010000001000110001";
wait for Clk_period;
Addr <= "0000001101010";
Trees_din <= "00000101000000000001010100000100";
wait for Clk_period;
Addr <= "0000001101011";
Trees_din <= "00000000000111100000001000110001";
wait for Clk_period;
Addr <= "0000001101100";
Trees_din <= "00000000000110000000001000110001";
wait for Clk_period;
Addr <= "0000001101101";
Trees_din <= "00000111000000000100010100100000";
wait for Clk_period;
Addr <= "0000001101110";
Trees_din <= "00000010000000000010010000010000";
wait for Clk_period;
Addr <= "0000001101111";
Trees_din <= "00000111000000000110000000001000";
wait for Clk_period;
Addr <= "0000001110000";
Trees_din <= "00000100000000000010100100000100";
wait for Clk_period;
Addr <= "0000001110001";
Trees_din <= "00000000010011010000001000110001";
wait for Clk_period;
Addr <= "0000001110010";
Trees_din <= "00000000001100010000001000110001";
wait for Clk_period;
Addr <= "0000001110011";
Trees_din <= "00000111000000000110001000000100";
wait for Clk_period;
Addr <= "0000001110100";
Trees_din <= "00000000010011110000001000110001";
wait for Clk_period;
Addr <= "0000001110101";
Trees_din <= "00000000001000010000001000110001";
wait for Clk_period;
Addr <= "0000001110110";
Trees_din <= "00000101000000000001000100001000";
wait for Clk_period;
Addr <= "0000001110111";
Trees_din <= "00000111000000000001101100000100";
wait for Clk_period;
Addr <= "0000001111000";
Trees_din <= "00000000001010000000001000110001";
wait for Clk_period;
Addr <= "0000001111001";
Trees_din <= "00000000000100010000001000110001";
wait for Clk_period;
Addr <= "0000001111010";
Trees_din <= "00000110000000000110001000000100";
wait for Clk_period;
Addr <= "0000001111011";
Trees_din <= "00000000011000000000001000110001";
wait for Clk_period;
Addr <= "0000001111100";
Trees_din <= "00000000001111100000001000110001";
wait for Clk_period;
Addr <= "0000001111101";
Trees_din <= "00000010000000000100010100010000";
wait for Clk_period;
Addr <= "0000001111110";
Trees_din <= "00000100000000000010101100001000";
wait for Clk_period;
Addr <= "0000001111111";
Trees_din <= "00000000000000000101001000000100";
wait for Clk_period;
Addr <= "0000010000000";
Trees_din <= "00000000000000000000001000110001";
wait for Clk_period;
Addr <= "0000010000001";
Trees_din <= "00000000010010110000001000110001";
wait for Clk_period;
Addr <= "0000010000010";
Trees_din <= "00000111000000000101010000000100";
wait for Clk_period;
Addr <= "0000010000011";
Trees_din <= "00000000000110000000001000110001";
wait for Clk_period;
Addr <= "0000010000100";
Trees_din <= "00000000010010100000001000110001";
wait for Clk_period;
Addr <= "0000010000101";
Trees_din <= "00000010000000000100001000001000";
wait for Clk_period;
Addr <= "0000010000110";
Trees_din <= "00000110000000000100000100000100";
wait for Clk_period;
Addr <= "0000010000111";
Trees_din <= "00000000000101010000001000110001";
wait for Clk_period;
Addr <= "0000010001000";
Trees_din <= "00000000000001000000001000110001";
wait for Clk_period;
Addr <= "0000010001001";
Trees_din <= "00000100000000000100000100000100";
wait for Clk_period;
Addr <= "0000010001010";
Trees_din <= "00000000001100110000001000110001";
wait for Clk_period;
Addr <= "0000010001011";
Trees_din <= "00000000001011110000001000110001";
wait for Clk_period;



----------tree 1-------------------

Addr <= "0000010001100";
Trees_din <= "00000111000000000000000010000000";
wait for Clk_period;
Addr <= "0000010001101";
Trees_din <= "00000110000000000000010001000000";
wait for Clk_period;
Addr <= "0000010001110";
Trees_din <= "00000011000000000000101000100000";
wait for Clk_period;
Addr <= "0000010001111";
Trees_din <= "00000001000000000101010100010000";
wait for Clk_period;
Addr <= "0000010010000";
Trees_din <= "00000110000000000011011000001000";
wait for Clk_period;
Addr <= "0000010010001";
Trees_din <= "00000111000000000011001000000100";
wait for Clk_period;
Addr <= "0000010010010";
Trees_din <= "00000000000001010000010000101111";
wait for Clk_period;
Addr <= "0000010010011";
Trees_din <= "00000000001110000000010000101111";
wait for Clk_period;
Addr <= "0000010010100";
Trees_din <= "00000110000000000101101100000100";
wait for Clk_period;
Addr <= "0000010010101";
Trees_din <= "00000000010100000000010000101111";
wait for Clk_period;
Addr <= "0000010010110";
Trees_din <= "00000000001111100000010000101111";
wait for Clk_period;
Addr <= "0000010010111";
Trees_din <= "00000101000000000010010100001000";
wait for Clk_period;
Addr <= "0000010011000";
Trees_din <= "00000000000000000000001000000100";
wait for Clk_period;
Addr <= "0000010011001";
Trees_din <= "00000000001001110000010000101111";
wait for Clk_period;
Addr <= "0000010011010";
Trees_din <= "00000000000110110000010000101111";
wait for Clk_period;
Addr <= "0000010011011";
Trees_din <= "00000001000000000000000100000100";
wait for Clk_period;
Addr <= "0000010011100";
Trees_din <= "00000000010101010000010000101111";
wait for Clk_period;
Addr <= "0000010011101";
Trees_din <= "00000000010001010000010000101111";
wait for Clk_period;
Addr <= "0000010011110";
Trees_din <= "00000010000000000110010000010000";
wait for Clk_period;
Addr <= "0000010011111";
Trees_din <= "00000001000000000101101100001000";
wait for Clk_period;
Addr <= "0000010100000";
Trees_din <= "00000011000000000011011100000100";
wait for Clk_period;
Addr <= "0000010100001";
Trees_din <= "00000000010111110000010000101111";
wait for Clk_period;
Addr <= "0000010100010";
Trees_din <= "00000000000101000000010000101111";
wait for Clk_period;
Addr <= "0000010100011";
Trees_din <= "00000010000000000011101000000100";
wait for Clk_period;
Addr <= "0000010100100";
Trees_din <= "00000000000110000000010000101111";
wait for Clk_period;
Addr <= "0000010100101";
Trees_din <= "00000000010010100000010000101111";
wait for Clk_period;
Addr <= "0000010100110";
Trees_din <= "00000111000000000101011100001000";
wait for Clk_period;
Addr <= "0000010100111";
Trees_din <= "00000000000000000010010100000100";
wait for Clk_period;
Addr <= "0000010101000";
Trees_din <= "00000000000111110000010000101111";
wait for Clk_period;
Addr <= "0000010101001";
Trees_din <= "00000000001111100000010000101111";
wait for Clk_period;
Addr <= "0000010101010";
Trees_din <= "00000000000000000000100000000100";
wait for Clk_period;
Addr <= "0000010101011";
Trees_din <= "00000000011001000000010000101111";
wait for Clk_period;
Addr <= "0000010101100";
Trees_din <= "00000000001111110000010000101111";
wait for Clk_period;
Addr <= "0000010101101";
Trees_din <= "00000001000000000110010000100000";
wait for Clk_period;
Addr <= "0000010101110";
Trees_din <= "00000100000000000101001000010000";
wait for Clk_period;
Addr <= "0000010101111";
Trees_din <= "00000111000000000000110100001000";
wait for Clk_period;
Addr <= "0000010110000";
Trees_din <= "00000111000000000010011000000100";
wait for Clk_period;
Addr <= "0000010110001";
Trees_din <= "00000000010100010000010000101111";
wait for Clk_period;
Addr <= "0000010110010";
Trees_din <= "00000000010010000000010000101111";
wait for Clk_period;
Addr <= "0000010110011";
Trees_din <= "00000010000000000100001100000100";
wait for Clk_period;
Addr <= "0000010110100";
Trees_din <= "00000000010011100000010000101111";
wait for Clk_period;
Addr <= "0000010110101";
Trees_din <= "00000000001100110000010000101111";
wait for Clk_period;
Addr <= "0000010110110";
Trees_din <= "00000001000000000100100100001000";
wait for Clk_period;
Addr <= "0000010110111";
Trees_din <= "00000111000000000010111100000100";
wait for Clk_period;
Addr <= "0000010111000";
Trees_din <= "00000000001011110000010000101111";
wait for Clk_period;
Addr <= "0000010111001";
Trees_din <= "00000000000000100000010000101111";
wait for Clk_period;
Addr <= "0000010111010";
Trees_din <= "00000110000000000001010100000100";
wait for Clk_period;
Addr <= "0000010111011";
Trees_din <= "00000000000111000000010000101111";
wait for Clk_period;
Addr <= "0000010111100";
Trees_din <= "00000000000000100000010000101111";
wait for Clk_period;
Addr <= "0000010111101";
Trees_din <= "00000011000000000000000000010000";
wait for Clk_period;
Addr <= "0000010111110";
Trees_din <= "00000110000000000100001100001000";
wait for Clk_period;
Addr <= "0000010111111";
Trees_din <= "00000000000000000010000100000100";
wait for Clk_period;
Addr <= "0000011000000";
Trees_din <= "00000000000111110000010000101111";
wait for Clk_period;
Addr <= "0000011000001";
Trees_din <= "00000000000000100000010000101111";
wait for Clk_period;
Addr <= "0000011000010";
Trees_din <= "00000000000000000101111100000100";
wait for Clk_period;
Addr <= "0000011000011";
Trees_din <= "00000000001001010000010000101111";
wait for Clk_period;
Addr <= "0000011000100";
Trees_din <= "00000000001100110000010000101111";
wait for Clk_period;
Addr <= "0000011000101";
Trees_din <= "00000011000000000001101000001000";
wait for Clk_period;
Addr <= "0000011000110";
Trees_din <= "00000101000000000011110000000100";
wait for Clk_period;
Addr <= "0000011000111";
Trees_din <= "00000000000100100000010000101111";
wait for Clk_period;
Addr <= "0000011001000";
Trees_din <= "00000000001010100000010000101111";
wait for Clk_period;
Addr <= "0000011001001";
Trees_din <= "00000111000000000101100100000100";
wait for Clk_period;
Addr <= "0000011001010";
Trees_din <= "00000000000111010000010000101111";
wait for Clk_period;
Addr <= "0000011001011";
Trees_din <= "00000000010001010000010000101111";
wait for Clk_period;
Addr <= "0000011001100";
Trees_din <= "00000111000000000010000101000000";
wait for Clk_period;
Addr <= "0000011001101";
Trees_din <= "00000100000000000000010000100000";
wait for Clk_period;
Addr <= "0000011001110";
Trees_din <= "00000110000000000000100000010000";
wait for Clk_period;
Addr <= "0000011001111";
Trees_din <= "00000001000000000000011100001000";
wait for Clk_period;
Addr <= "0000011010000";
Trees_din <= "00000111000000000010000000000100";
wait for Clk_period;
Addr <= "0000011010001";
Trees_din <= "00000000010111000000010000101111";
wait for Clk_period;
Addr <= "0000011010010";
Trees_din <= "00000000010010010000010000101111";
wait for Clk_period;
Addr <= "0000011010011";
Trees_din <= "00000000000000000011010100000100";
wait for Clk_period;
Addr <= "0000011010100";
Trees_din <= "00000000001110000000010000101111";
wait for Clk_period;
Addr <= "0000011010101";
Trees_din <= "00000000001101110000010000101111";
wait for Clk_period;
Addr <= "0000011010110";
Trees_din <= "00000111000000000011100000001000";
wait for Clk_period;
Addr <= "0000011010111";
Trees_din <= "00000101000000000011011100000100";
wait for Clk_period;
Addr <= "0000011011000";
Trees_din <= "00000000000000100000010000101111";
wait for Clk_period;
Addr <= "0000011011001";
Trees_din <= "00000000000010000000010000101111";
wait for Clk_period;
Addr <= "0000011011010";
Trees_din <= "00000001000000000101001000000100";
wait for Clk_period;
Addr <= "0000011011011";
Trees_din <= "00000000001111110000010000101111";
wait for Clk_period;
Addr <= "0000011011100";
Trees_din <= "00000000001010110000010000101111";
wait for Clk_period;
Addr <= "0000011011101";
Trees_din <= "00000100000000000001110000010000";
wait for Clk_period;
Addr <= "0000011011110";
Trees_din <= "00000000000000000001001000001000";
wait for Clk_period;
Addr <= "0000011011111";
Trees_din <= "00000101000000000100000000000100";
wait for Clk_period;
Addr <= "0000011100000";
Trees_din <= "00000000001000010000010000101111";
wait for Clk_period;
Addr <= "0000011100001";
Trees_din <= "00000000000010000000010000101111";
wait for Clk_period;
Addr <= "0000011100010";
Trees_din <= "00000001000000000100100000000100";
wait for Clk_period;
Addr <= "0000011100011";
Trees_din <= "00000000001110000000010000101111";
wait for Clk_period;
Addr <= "0000011100100";
Trees_din <= "00000000001100010000010000101111";
wait for Clk_period;
Addr <= "0000011100101";
Trees_din <= "00000101000000000110001000001000";
wait for Clk_period;
Addr <= "0000011100110";
Trees_din <= "00000111000000000010110000000100";
wait for Clk_period;
Addr <= "0000011100111";
Trees_din <= "00000000001111100000010000101111";
wait for Clk_period;
Addr <= "0000011101000";
Trees_din <= "00000000010011010000010000101111";
wait for Clk_period;
Addr <= "0000011101001";
Trees_din <= "00000001000000000010010000000100";
wait for Clk_period;
Addr <= "0000011101010";
Trees_din <= "00000000001100110000010000101111";
wait for Clk_period;
Addr <= "0000011101011";
Trees_din <= "00000000001011000000010000101111";
wait for Clk_period;
Addr <= "0000011101100";
Trees_din <= "00000101000000000011001100100000";
wait for Clk_period;
Addr <= "0000011101101";
Trees_din <= "00000100000000000010100100010000";
wait for Clk_period;
Addr <= "0000011101110";
Trees_din <= "00000110000000000001100000001000";
wait for Clk_period;
Addr <= "0000011101111";
Trees_din <= "00000001000000000000110100000100";
wait for Clk_period;
Addr <= "0000011110000";
Trees_din <= "00000000000111000000010000101111";
wait for Clk_period;
Addr <= "0000011110001";
Trees_din <= "00000000001011110000010000101111";
wait for Clk_period;
Addr <= "0000011110010";
Trees_din <= "00000111000000000011010000000100";
wait for Clk_period;
Addr <= "0000011110011";
Trees_din <= "00000000001110100000010000101111";
wait for Clk_period;
Addr <= "0000011110100";
Trees_din <= "00000000010000010000010000101111";
wait for Clk_period;
Addr <= "0000011110101";
Trees_din <= "00000001000000000100011000001000";
wait for Clk_period;
Addr <= "0000011110110";
Trees_din <= "00000100000000000010100000000100";
wait for Clk_period;
Addr <= "0000011110111";
Trees_din <= "00000000001100110000010000101111";
wait for Clk_period;
Addr <= "0000011111000";
Trees_din <= "00000000001100000000010000101111";
wait for Clk_period;
Addr <= "0000011111001";
Trees_din <= "00000000000000000000001100000100";
wait for Clk_period;
Addr <= "0000011111010";
Trees_din <= "00000000010000010000010000101111";
wait for Clk_period;
Addr <= "0000011111011";
Trees_din <= "00000000000100010000010000101111";
wait for Clk_period;
Addr <= "0000011111100";
Trees_din <= "00000000000000000000000100010000";
wait for Clk_period;
Addr <= "0000011111101";
Trees_din <= "00000110000000000100011000001000";
wait for Clk_period;
Addr <= "0000011111110";
Trees_din <= "00000111000000000010001100000100";
wait for Clk_period;
Addr <= "0000011111111";
Trees_din <= "00000000001001010000010000101111";
wait for Clk_period;
Addr <= "0000100000000";
Trees_din <= "00000000000000010000010000101111";
wait for Clk_period;
Addr <= "0000100000001";
Trees_din <= "00000101000000000001100000000100";
wait for Clk_period;
Addr <= "0000100000010";
Trees_din <= "00000000010101110000010000101111";
wait for Clk_period;
Addr <= "0000100000011";
Trees_din <= "00000000001001010000010000101111";
wait for Clk_period;
Addr <= "0000100000100";
Trees_din <= "00000001000000000000001100001000";
wait for Clk_period;
Addr <= "0000100000101";
Trees_din <= "00000101000000000100011000000100";
wait for Clk_period;
Addr <= "0000100000110";
Trees_din <= "00000000001000110000010000101111";
wait for Clk_period;
Addr <= "0000100000111";
Trees_din <= "00000000000111100000010000101111";
wait for Clk_period;
Addr <= "0000100001000";
Trees_din <= "00000010000000000000010100000100";
wait for Clk_period;
Addr <= "0000100001001";
Trees_din <= "00000000001101100000010000101111";
wait for Clk_period;
Addr <= "0000100001010";
Trees_din <= "00000000001110010000010000101111";
wait for Clk_period;



----------tree 2-------------------

Addr <= "0000100001011";
Trees_din <= "00000101000000000010101110000000";
wait for Clk_period;
Addr <= "0000100001100";
Trees_din <= "00000011000000000001011001000000";
wait for Clk_period;
Addr <= "0000100001101";
Trees_din <= "00000000000000000100101100100000";
wait for Clk_period;
Addr <= "0000100001110";
Trees_din <= "00000110000000000001011000010000";
wait for Clk_period;
Addr <= "0000100001111";
Trees_din <= "00000000000000000010001000001000";
wait for Clk_period;
Addr <= "0000100010000";
Trees_din <= "00000100000000000011110100000100";
wait for Clk_period;
Addr <= "0000100010001";
Trees_din <= "00000000001110110000011000101001";
wait for Clk_period;
Addr <= "0000100010010";
Trees_din <= "00000000001011010000011000101001";
wait for Clk_period;
Addr <= "0000100010011";
Trees_din <= "00000110000000000100110000000100";
wait for Clk_period;
Addr <= "0000100010100";
Trees_din <= "00000000010110110000011000101001";
wait for Clk_period;
Addr <= "0000100010101";
Trees_din <= "00000000001101100000011000101001";
wait for Clk_period;
Addr <= "0000100010110";
Trees_din <= "00000111000000000100100100001000";
wait for Clk_period;
Addr <= "0000100010111";
Trees_din <= "00000110000000000110001000000100";
wait for Clk_period;
Addr <= "0000100011000";
Trees_din <= "00000000000000010000011000101001";
wait for Clk_period;
Addr <= "0000100011001";
Trees_din <= "00000000000011110000011000101001";
wait for Clk_period;
Addr <= "0000100011010";
Trees_din <= "00000001000000000101101000000100";
wait for Clk_period;
Addr <= "0000100011011";
Trees_din <= "00000000001011110000011000101001";
wait for Clk_period;
Addr <= "0000100011100";
Trees_din <= "00000000000000110000011000101001";
wait for Clk_period;
Addr <= "0000100011101";
Trees_din <= "00000110000000000001101100010000";
wait for Clk_period;
Addr <= "0000100011110";
Trees_din <= "00000110000000000101100000001000";
wait for Clk_period;
Addr <= "0000100011111";
Trees_din <= "00000101000000000100100100000100";
wait for Clk_period;
Addr <= "0000100100000";
Trees_din <= "00000000001001000000011000101001";
wait for Clk_period;
Addr <= "0000100100001";
Trees_din <= "00000000010110100000011000101001";
wait for Clk_period;
Addr <= "0000100100010";
Trees_din <= "00000111000000000100110100000100";
wait for Clk_period;
Addr <= "0000100100011";
Trees_din <= "00000000000011110000011000101001";
wait for Clk_period;
Addr <= "0000100100100";
Trees_din <= "00000000010110000000011000101001";
wait for Clk_period;
Addr <= "0000100100101";
Trees_din <= "00000101000000000001011100001000";
wait for Clk_period;
Addr <= "0000100100110";
Trees_din <= "00000001000000000110001000000100";
wait for Clk_period;
Addr <= "0000100100111";
Trees_din <= "00000000001101000000011000101001";
wait for Clk_period;
Addr <= "0000100101000";
Trees_din <= "00000000000010110000011000101001";
wait for Clk_period;
Addr <= "0000100101001";
Trees_din <= "00000001000000000000111100000100";
wait for Clk_period;
Addr <= "0000100101010";
Trees_din <= "00000000001001000000011000101001";
wait for Clk_period;
Addr <= "0000100101011";
Trees_din <= "00000000010100110000011000101001";
wait for Clk_period;
Addr <= "0000100101100";
Trees_din <= "00000110000000000011001000100000";
wait for Clk_period;
Addr <= "0000100101101";
Trees_din <= "00000010000000000101101100010000";
wait for Clk_period;
Addr <= "0000100101110";
Trees_din <= "00000111000000000100001100001000";
wait for Clk_period;
Addr <= "0000100101111";
Trees_din <= "00000101000000000100000100000100";
wait for Clk_period;
Addr <= "0000100110000";
Trees_din <= "00000000001100010000011000101001";
wait for Clk_period;
Addr <= "0000100110001";
Trees_din <= "00000000000111000000011000101001";
wait for Clk_period;
Addr <= "0000100110010";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "0000100110011";
Trees_din <= "00000000000101000000011000101001";
wait for Clk_period;
Addr <= "0000100110100";
Trees_din <= "00000000000101110000011000101001";
wait for Clk_period;
Addr <= "0000100110101";
Trees_din <= "00000010000000000101101000001000";
wait for Clk_period;
Addr <= "0000100110110";
Trees_din <= "00000001000000000110000100000100";
wait for Clk_period;
Addr <= "0000100110111";
Trees_din <= "00000000000111010000011000101001";
wait for Clk_period;
Addr <= "0000100111000";
Trees_din <= "00000000000001010000011000101001";
wait for Clk_period;
Addr <= "0000100111001";
Trees_din <= "00000100000000000011011100000100";
wait for Clk_period;
Addr <= "0000100111010";
Trees_din <= "00000000001011000000011000101001";
wait for Clk_period;
Addr <= "0000100111011";
Trees_din <= "00000000010010100000011000101001";
wait for Clk_period;
Addr <= "0000100111100";
Trees_din <= "00000111000000000000111000010000";
wait for Clk_period;
Addr <= "0000100111101";
Trees_din <= "00000111000000000000001000001000";
wait for Clk_period;
Addr <= "0000100111110";
Trees_din <= "00000010000000000011011100000100";
wait for Clk_period;
Addr <= "0000100111111";
Trees_din <= "00000000000000000000011000101001";
wait for Clk_period;
Addr <= "0000101000000";
Trees_din <= "00000000000000110000011000101001";
wait for Clk_period;
Addr <= "0000101000001";
Trees_din <= "00000010000000000100101100000100";
wait for Clk_period;
Addr <= "0000101000010";
Trees_din <= "00000000010100010000011000101001";
wait for Clk_period;
Addr <= "0000101000011";
Trees_din <= "00000000010110110000011000101001";
wait for Clk_period;
Addr <= "0000101000100";
Trees_din <= "00000111000000000000110000001000";
wait for Clk_period;
Addr <= "0000101000101";
Trees_din <= "00000100000000000000110100000100";
wait for Clk_period;
Addr <= "0000101000110";
Trees_din <= "00000000001111110000011000101001";
wait for Clk_period;
Addr <= "0000101000111";
Trees_din <= "00000000000100110000011000101001";
wait for Clk_period;
Addr <= "0000101001000";
Trees_din <= "00000001000000000000001100000100";
wait for Clk_period;
Addr <= "0000101001001";
Trees_din <= "00000000010000100000011000101001";
wait for Clk_period;
Addr <= "0000101001010";
Trees_din <= "00000000000110100000011000101001";
wait for Clk_period;
Addr <= "0000101001011";
Trees_din <= "00000000000000000000110101000000";
wait for Clk_period;
Addr <= "0000101001100";
Trees_din <= "00000100000000000010001000100000";
wait for Clk_period;
Addr <= "0000101001101";
Trees_din <= "00000010000000000100001000010000";
wait for Clk_period;
Addr <= "0000101001110";
Trees_din <= "00000001000000000100100000001000";
wait for Clk_period;
Addr <= "0000101001111";
Trees_din <= "00000011000000000000001000000100";
wait for Clk_period;
Addr <= "0000101010000";
Trees_din <= "00000000010111100000011000101001";
wait for Clk_period;
Addr <= "0000101010001";
Trees_din <= "00000000000010110000011000101001";
wait for Clk_period;
Addr <= "0000101010010";
Trees_din <= "00000111000000000001000000000100";
wait for Clk_period;
Addr <= "0000101010011";
Trees_din <= "00000000000000010000011000101001";
wait for Clk_period;
Addr <= "0000101010100";
Trees_din <= "00000000001010110000011000101001";
wait for Clk_period;
Addr <= "0000101010101";
Trees_din <= "00000011000000000100010100001000";
wait for Clk_period;
Addr <= "0000101010110";
Trees_din <= "00000110000000000011000100000100";
wait for Clk_period;
Addr <= "0000101010111";
Trees_din <= "00000000010111000000011000101001";
wait for Clk_period;
Addr <= "0000101011000";
Trees_din <= "00000000010010110000011000101001";
wait for Clk_period;
Addr <= "0000101011001";
Trees_din <= "00000111000000000010110000000100";
wait for Clk_period;
Addr <= "0000101011010";
Trees_din <= "00000000001011110000011000101001";
wait for Clk_period;
Addr <= "0000101011011";
Trees_din <= "00000000001001010000011000101001";
wait for Clk_period;
Addr <= "0000101011100";
Trees_din <= "00000010000000000110001000010000";
wait for Clk_period;
Addr <= "0000101011101";
Trees_din <= "00000010000000000000100100001000";
wait for Clk_period;
Addr <= "0000101011110";
Trees_din <= "00000000000000000101100100000100";
wait for Clk_period;
Addr <= "0000101011111";
Trees_din <= "00000000010001000000011000101001";
wait for Clk_period;
Addr <= "0000101100000";
Trees_din <= "00000000001001100000011000101001";
wait for Clk_period;
Addr <= "0000101100001";
Trees_din <= "00000010000000000101011100000100";
wait for Clk_period;
Addr <= "0000101100010";
Trees_din <= "00000000010010000000011000101001";
wait for Clk_period;
Addr <= "0000101100011";
Trees_din <= "00000000010011000000011000101001";
wait for Clk_period;
Addr <= "0000101100100";
Trees_din <= "00000000000000000011000100001000";
wait for Clk_period;
Addr <= "0000101100101";
Trees_din <= "00000101000000000011101100000100";
wait for Clk_period;
Addr <= "0000101100110";
Trees_din <= "00000000000001100000011000101001";
wait for Clk_period;
Addr <= "0000101100111";
Trees_din <= "00000000010101100000011000101001";
wait for Clk_period;
Addr <= "0000101101000";
Trees_din <= "00000110000000000001000000000100";
wait for Clk_period;
Addr <= "0000101101001";
Trees_din <= "00000000001110110000011000101001";
wait for Clk_period;
Addr <= "0000101101010";
Trees_din <= "00000000001111110000011000101001";
wait for Clk_period;
Addr <= "0000101101011";
Trees_din <= "00000000000000000010111000100000";
wait for Clk_period;
Addr <= "0000101101100";
Trees_din <= "00000110000000000000111100010000";
wait for Clk_period;
Addr <= "0000101101101";
Trees_din <= "00000010000000000101011100001000";
wait for Clk_period;
Addr <= "0000101101110";
Trees_din <= "00000010000000000101011100000100";
wait for Clk_period;
Addr <= "0000101101111";
Trees_din <= "00000000001001100000011000101001";
wait for Clk_period;
Addr <= "0000101110000";
Trees_din <= "00000000000100110000011000101001";
wait for Clk_period;
Addr <= "0000101110001";
Trees_din <= "00000100000000000101111100000100";
wait for Clk_period;
Addr <= "0000101110010";
Trees_din <= "00000000000001100000011000101001";
wait for Clk_period;
Addr <= "0000101110011";
Trees_din <= "00000000010101000000011000101001";
wait for Clk_period;
Addr <= "0000101110100";
Trees_din <= "00000110000000000011101000001000";
wait for Clk_period;
Addr <= "0000101110101";
Trees_din <= "00000111000000000101010000000100";
wait for Clk_period;
Addr <= "0000101110110";
Trees_din <= "00000000000010010000011000101001";
wait for Clk_period;
Addr <= "0000101110111";
Trees_din <= "00000000001110100000011000101001";
wait for Clk_period;
Addr <= "0000101111000";
Trees_din <= "00000101000000000101000000000100";
wait for Clk_period;
Addr <= "0000101111001";
Trees_din <= "00000000001110010000011000101001";
wait for Clk_period;
Addr <= "0000101111010";
Trees_din <= "00000000001111100000011000101001";
wait for Clk_period;
Addr <= "0000101111011";
Trees_din <= "00000001000000000100111100010000";
wait for Clk_period;
Addr <= "0000101111100";
Trees_din <= "00000011000000000100000000001000";
wait for Clk_period;
Addr <= "0000101111101";
Trees_din <= "00000010000000000001011000000100";
wait for Clk_period;
Addr <= "0000101111110";
Trees_din <= "00000000001100100000011000101001";
wait for Clk_period;
Addr <= "0000101111111";
Trees_din <= "00000000001110100000011000101001";
wait for Clk_period;
Addr <= "0000110000000";
Trees_din <= "00000110000000000010011100000100";
wait for Clk_period;
Addr <= "0000110000001";
Trees_din <= "00000000010000000000011000101001";
wait for Clk_period;
Addr <= "0000110000010";
Trees_din <= "00000000001010010000011000101001";
wait for Clk_period;
Addr <= "0000110000011";
Trees_din <= "00000010000000000100001100001000";
wait for Clk_period;
Addr <= "0000110000100";
Trees_din <= "00000100000000000001100000000100";
wait for Clk_period;
Addr <= "0000110000101";
Trees_din <= "00000000001111100000011000101001";
wait for Clk_period;
Addr <= "0000110000110";
Trees_din <= "00000000001111110000011000101001";
wait for Clk_period;
Addr <= "0000110000111";
Trees_din <= "00000001000000000001001100000100";
wait for Clk_period;
Addr <= "0000110001000";
Trees_din <= "00000000001101000000011000101001";
wait for Clk_period;
Addr <= "0000110001001";
Trees_din <= "00000000001000110000011000101001";
wait for Clk_period;



----------tree 3-------------------

Addr <= "0000110001010";
Trees_din <= "00000111000000000010001110000000";
wait for Clk_period;
Addr <= "0000110001011";
Trees_din <= "00000100000000000100100001000000";
wait for Clk_period;
Addr <= "0000110001100";
Trees_din <= "00000111000000000000101000100000";
wait for Clk_period;
Addr <= "0000110001101";
Trees_din <= "00000110000000000001000000010000";
wait for Clk_period;
Addr <= "0000110001110";
Trees_din <= "00000011000000000010110100001000";
wait for Clk_period;
Addr <= "0000110001111";
Trees_din <= "00000111000000000001110000000100";
wait for Clk_period;
Addr <= "0000110010000";
Trees_din <= "00000000001011010000100000100111";
wait for Clk_period;
Addr <= "0000110010001";
Trees_din <= "00000000010111110000100000100111";
wait for Clk_period;
Addr <= "0000110010010";
Trees_din <= "00000111000000000001010100000100";
wait for Clk_period;
Addr <= "0000110010011";
Trees_din <= "00000000001111010000100000100111";
wait for Clk_period;
Addr <= "0000110010100";
Trees_din <= "00000000010110110000100000100111";
wait for Clk_period;
Addr <= "0000110010101";
Trees_din <= "00000000000000000100001100001000";
wait for Clk_period;
Addr <= "0000110010110";
Trees_din <= "00000110000000000100010000000100";
wait for Clk_period;
Addr <= "0000110010111";
Trees_din <= "00000000010000100000100000100111";
wait for Clk_period;
Addr <= "0000110011000";
Trees_din <= "00000000001000000000100000100111";
wait for Clk_period;
Addr <= "0000110011001";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "0000110011010";
Trees_din <= "00000000010001100000100000100111";
wait for Clk_period;
Addr <= "0000110011011";
Trees_din <= "00000000010101110000100000100111";
wait for Clk_period;
Addr <= "0000110011100";
Trees_din <= "00000100000000000100001000010000";
wait for Clk_period;
Addr <= "0000110011101";
Trees_din <= "00000011000000000101111100001000";
wait for Clk_period;
Addr <= "0000110011110";
Trees_din <= "00000011000000000000101100000100";
wait for Clk_period;
Addr <= "0000110011111";
Trees_din <= "00000000010010000000100000100111";
wait for Clk_period;
Addr <= "0000110100000";
Trees_din <= "00000000000011110000100000100111";
wait for Clk_period;
Addr <= "0000110100001";
Trees_din <= "00000100000000000010001000000100";
wait for Clk_period;
Addr <= "0000110100010";
Trees_din <= "00000000010100110000100000100111";
wait for Clk_period;
Addr <= "0000110100011";
Trees_din <= "00000000010111110000100000100111";
wait for Clk_period;
Addr <= "0000110100100";
Trees_din <= "00000111000000000110001100001000";
wait for Clk_period;
Addr <= "0000110100101";
Trees_din <= "00000001000000000000000000000100";
wait for Clk_period;
Addr <= "0000110100110";
Trees_din <= "00000000000011000000100000100111";
wait for Clk_period;
Addr <= "0000110100111";
Trees_din <= "00000000000110010000100000100111";
wait for Clk_period;
Addr <= "0000110101000";
Trees_din <= "00000000000000000010101000000100";
wait for Clk_period;
Addr <= "0000110101001";
Trees_din <= "00000000001010000000100000100111";
wait for Clk_period;
Addr <= "0000110101010";
Trees_din <= "00000000001111000000100000100111";
wait for Clk_period;
Addr <= "0000110101011";
Trees_din <= "00000011000000000010001000100000";
wait for Clk_period;
Addr <= "0000110101100";
Trees_din <= "00000010000000000000000000010000";
wait for Clk_period;
Addr <= "0000110101101";
Trees_din <= "00000000000000000000100000001000";
wait for Clk_period;
Addr <= "0000110101110";
Trees_din <= "00000011000000000011010000000100";
wait for Clk_period;
Addr <= "0000110101111";
Trees_din <= "00000000000111100000100000100111";
wait for Clk_period;
Addr <= "0000110110000";
Trees_din <= "00000000010000010000100000100111";
wait for Clk_period;
Addr <= "0000110110001";
Trees_din <= "00000110000000000100101100000100";
wait for Clk_period;
Addr <= "0000110110010";
Trees_din <= "00000000001010010000100000100111";
wait for Clk_period;
Addr <= "0000110110011";
Trees_din <= "00000000010010000000100000100111";
wait for Clk_period;
Addr <= "0000110110100";
Trees_din <= "00000110000000000011010100001000";
wait for Clk_period;
Addr <= "0000110110101";
Trees_din <= "00000111000000000101000000000100";
wait for Clk_period;
Addr <= "0000110110110";
Trees_din <= "00000000010100010000100000100111";
wait for Clk_period;
Addr <= "0000110110111";
Trees_din <= "00000000011000000000100000100111";
wait for Clk_period;
Addr <= "0000110111000";
Trees_din <= "00000110000000000000100100000100";
wait for Clk_period;
Addr <= "0000110111001";
Trees_din <= "00000000001110010000100000100111";
wait for Clk_period;
Addr <= "0000110111010";
Trees_din <= "00000000000010110000100000100111";
wait for Clk_period;
Addr <= "0000110111011";
Trees_din <= "00000110000000000001111100010000";
wait for Clk_period;
Addr <= "0000110111100";
Trees_din <= "00000100000000000011111100001000";
wait for Clk_period;
Addr <= "0000110111101";
Trees_din <= "00000111000000000100001000000100";
wait for Clk_period;
Addr <= "0000110111110";
Trees_din <= "00000000010011110000100000100111";
wait for Clk_period;
Addr <= "0000110111111";
Trees_din <= "00000000000100000000100000100111";
wait for Clk_period;
Addr <= "0000111000000";
Trees_din <= "00000001000000000011110000000100";
wait for Clk_period;
Addr <= "0000111000001";
Trees_din <= "00000000000001100000100000100111";
wait for Clk_period;
Addr <= "0000111000010";
Trees_din <= "00000000001001100000100000100111";
wait for Clk_period;
Addr <= "0000111000011";
Trees_din <= "00000001000000000000001000001000";
wait for Clk_period;
Addr <= "0000111000100";
Trees_din <= "00000110000000000010111000000100";
wait for Clk_period;
Addr <= "0000111000101";
Trees_din <= "00000000001111100000100000100111";
wait for Clk_period;
Addr <= "0000111000110";
Trees_din <= "00000000000000110000100000100111";
wait for Clk_period;
Addr <= "0000111000111";
Trees_din <= "00000100000000000010011000000100";
wait for Clk_period;
Addr <= "0000111001000";
Trees_din <= "00000000000000100000100000100111";
wait for Clk_period;
Addr <= "0000111001001";
Trees_din <= "00000000001011100000100000100111";
wait for Clk_period;
Addr <= "0000111001010";
Trees_din <= "00000000000000000000010101000000";
wait for Clk_period;
Addr <= "0000111001011";
Trees_din <= "00000110000000000100100100100000";
wait for Clk_period;
Addr <= "0000111001100";
Trees_din <= "00000111000000000010001100010000";
wait for Clk_period;
Addr <= "0000111001101";
Trees_din <= "00000011000000000101010000001000";
wait for Clk_period;
Addr <= "0000111001110";
Trees_din <= "00000011000000000010110000000100";
wait for Clk_period;
Addr <= "0000111001111";
Trees_din <= "00000000000101100000100000100111";
wait for Clk_period;
Addr <= "0000111010000";
Trees_din <= "00000000010100100000100000100111";
wait for Clk_period;
Addr <= "0000111010001";
Trees_din <= "00000001000000000011110100000100";
wait for Clk_period;
Addr <= "0000111010010";
Trees_din <= "00000000001001010000100000100111";
wait for Clk_period;
Addr <= "0000111010011";
Trees_din <= "00000000010000010000100000100111";
wait for Clk_period;
Addr <= "0000111010100";
Trees_din <= "00000000000000000110001100001000";
wait for Clk_period;
Addr <= "0000111010101";
Trees_din <= "00000100000000000001001000000100";
wait for Clk_period;
Addr <= "0000111010110";
Trees_din <= "00000000011001000000100000100111";
wait for Clk_period;
Addr <= "0000111010111";
Trees_din <= "00000000010011100000100000100111";
wait for Clk_period;
Addr <= "0000111011000";
Trees_din <= "00000100000000000001101000000100";
wait for Clk_period;
Addr <= "0000111011001";
Trees_din <= "00000000001000010000100000100111";
wait for Clk_period;
Addr <= "0000111011010";
Trees_din <= "00000000000001110000100000100111";
wait for Clk_period;
Addr <= "0000111011011";
Trees_din <= "00000111000000000000000100010000";
wait for Clk_period;
Addr <= "0000111011100";
Trees_din <= "00000100000000000101111000001000";
wait for Clk_period;
Addr <= "0000111011101";
Trees_din <= "00000001000000000101010000000100";
wait for Clk_period;
Addr <= "0000111011110";
Trees_din <= "00000000010001010000100000100111";
wait for Clk_period;
Addr <= "0000111011111";
Trees_din <= "00000000010010100000100000100111";
wait for Clk_period;
Addr <= "0000111100000";
Trees_din <= "00000110000000000101100100000100";
wait for Clk_period;
Addr <= "0000111100001";
Trees_din <= "00000000000100000000100000100111";
wait for Clk_period;
Addr <= "0000111100010";
Trees_din <= "00000000000001110000100000100111";
wait for Clk_period;
Addr <= "0000111100011";
Trees_din <= "00000100000000000001001000001000";
wait for Clk_period;
Addr <= "0000111100100";
Trees_din <= "00000111000000000011010000000100";
wait for Clk_period;
Addr <= "0000111100101";
Trees_din <= "00000000000101000000100000100111";
wait for Clk_period;
Addr <= "0000111100110";
Trees_din <= "00000000000110010000100000100111";
wait for Clk_period;
Addr <= "0000111100111";
Trees_din <= "00000000000000000101110000000100";
wait for Clk_period;
Addr <= "0000111101000";
Trees_din <= "00000000000001000000100000100111";
wait for Clk_period;
Addr <= "0000111101001";
Trees_din <= "00000000000111010000100000100111";
wait for Clk_period;
Addr <= "0000111101010";
Trees_din <= "00000111000000000000100100100000";
wait for Clk_period;
Addr <= "0000111101011";
Trees_din <= "00000101000000000000011100010000";
wait for Clk_period;
Addr <= "0000111101100";
Trees_din <= "00000000000000000000101100001000";
wait for Clk_period;
Addr <= "0000111101101";
Trees_din <= "00000110000000000000101100000100";
wait for Clk_period;
Addr <= "0000111101110";
Trees_din <= "00000000010010100000100000100111";
wait for Clk_period;
Addr <= "0000111101111";
Trees_din <= "00000000010001000000100000100111";
wait for Clk_period;
Addr <= "0000111110000";
Trees_din <= "00000000000000000000000100000100";
wait for Clk_period;
Addr <= "0000111110001";
Trees_din <= "00000000010101000000100000100111";
wait for Clk_period;
Addr <= "0000111110010";
Trees_din <= "00000000000100010000100000100111";
wait for Clk_period;
Addr <= "0000111110011";
Trees_din <= "00000001000000000000001000001000";
wait for Clk_period;
Addr <= "0000111110100";
Trees_din <= "00000010000000000011001000000100";
wait for Clk_period;
Addr <= "0000111110101";
Trees_din <= "00000000000111110000100000100111";
wait for Clk_period;
Addr <= "0000111110110";
Trees_din <= "00000000010111010000100000100111";
wait for Clk_period;
Addr <= "0000111110111";
Trees_din <= "00000100000000000011001000000100";
wait for Clk_period;
Addr <= "0000111111000";
Trees_din <= "00000000000000100000100000100111";
wait for Clk_period;
Addr <= "0000111111001";
Trees_din <= "00000000001101110000100000100111";
wait for Clk_period;
Addr <= "0000111111010";
Trees_din <= "00000100000000000101010000010000";
wait for Clk_period;
Addr <= "0000111111011";
Trees_din <= "00000000000000000101010100001000";
wait for Clk_period;
Addr <= "0000111111100";
Trees_din <= "00000110000000000011001100000100";
wait for Clk_period;
Addr <= "0000111111101";
Trees_din <= "00000000010101110000100000100111";
wait for Clk_period;
Addr <= "0000111111110";
Trees_din <= "00000000010101110000100000100111";
wait for Clk_period;
Addr <= "0000111111111";
Trees_din <= "00000011000000000100110100000100";
wait for Clk_period;
Addr <= "0001000000000";
Trees_din <= "00000000000100110000100000100111";
wait for Clk_period;
Addr <= "0001000000001";
Trees_din <= "00000000000111000000100000100111";
wait for Clk_period;
Addr <= "0001000000010";
Trees_din <= "00000100000000000001001100001000";
wait for Clk_period;
Addr <= "0001000000011";
Trees_din <= "00000111000000000011101000000100";
wait for Clk_period;
Addr <= "0001000000100";
Trees_din <= "00000000001101110000100000100111";
wait for Clk_period;
Addr <= "0001000000101";
Trees_din <= "00000000001110100000100000100111";
wait for Clk_period;
Addr <= "0001000000110";
Trees_din <= "00000110000000000001010000000100";
wait for Clk_period;
Addr <= "0001000000111";
Trees_din <= "00000000010011110000100000100111";
wait for Clk_period;
Addr <= "0001000001000";
Trees_din <= "00000000001101100000100000100111";
wait for Clk_period;



----------tree 4-------------------

Addr <= "0001000001001";
Trees_din <= "00000111000000000100101010000000";
wait for Clk_period;
Addr <= "0001000001010";
Trees_din <= "00000100000000000001010001000000";
wait for Clk_period;
Addr <= "0001000001011";
Trees_din <= "00000111000000000110001000100000";
wait for Clk_period;
Addr <= "0001000001100";
Trees_din <= "00000110000000000100101100010000";
wait for Clk_period;
Addr <= "0001000001101";
Trees_din <= "00000000000000000110001100001000";
wait for Clk_period;
Addr <= "0001000001110";
Trees_din <= "00000111000000000000101000000100";
wait for Clk_period;
Addr <= "0001000001111";
Trees_din <= "00000000011000010000101000100001";
wait for Clk_period;
Addr <= "0001000010000";
Trees_din <= "00000000010010010000101000100001";
wait for Clk_period;
Addr <= "0001000010001";
Trees_din <= "00000000000000000100001100000100";
wait for Clk_period;
Addr <= "0001000010010";
Trees_din <= "00000000000100110000101000100001";
wait for Clk_period;
Addr <= "0001000010011";
Trees_din <= "00000000000101110000101000100001";
wait for Clk_period;
Addr <= "0001000010100";
Trees_din <= "00000000000000000011100000001000";
wait for Clk_period;
Addr <= "0001000010101";
Trees_din <= "00000110000000000101100000000100";
wait for Clk_period;
Addr <= "0001000010110";
Trees_din <= "00000000010001110000101000100001";
wait for Clk_period;
Addr <= "0001000010111";
Trees_din <= "00000000001100100000101000100001";
wait for Clk_period;
Addr <= "0001000011000";
Trees_din <= "00000010000000000011011100000100";
wait for Clk_period;
Addr <= "0001000011001";
Trees_din <= "00000000001111000000101000100001";
wait for Clk_period;
Addr <= "0001000011010";
Trees_din <= "00000000001010100000101000100001";
wait for Clk_period;
Addr <= "0001000011011";
Trees_din <= "00000000000000000011001100010000";
wait for Clk_period;
Addr <= "0001000011100";
Trees_din <= "00000100000000000100011000001000";
wait for Clk_period;
Addr <= "0001000011101";
Trees_din <= "00000001000000000000100100000100";
wait for Clk_period;
Addr <= "0001000011110";
Trees_din <= "00000000010000000000101000100001";
wait for Clk_period;
Addr <= "0001000011111";
Trees_din <= "00000000010011100000101000100001";
wait for Clk_period;
Addr <= "0001000100000";
Trees_din <= "00000110000000000001100000000100";
wait for Clk_period;
Addr <= "0001000100001";
Trees_din <= "00000000001110100000101000100001";
wait for Clk_period;
Addr <= "0001000100010";
Trees_din <= "00000000001110010000101000100001";
wait for Clk_period;
Addr <= "0001000100011";
Trees_din <= "00000100000000000010111000001000";
wait for Clk_period;
Addr <= "0001000100100";
Trees_din <= "00000100000000000101001100000100";
wait for Clk_period;
Addr <= "0001000100101";
Trees_din <= "00000000000011100000101000100001";
wait for Clk_period;
Addr <= "0001000100110";
Trees_din <= "00000000000010100000101000100001";
wait for Clk_period;
Addr <= "0001000100111";
Trees_din <= "00000100000000000011000100000100";
wait for Clk_period;
Addr <= "0001000101000";
Trees_din <= "00000000011001000000101000100001";
wait for Clk_period;
Addr <= "0001000101001";
Trees_din <= "00000000010100100000101000100001";
wait for Clk_period;
Addr <= "0001000101010";
Trees_din <= "00000101000000000011110000100000";
wait for Clk_period;
Addr <= "0001000101011";
Trees_din <= "00000000000000000101010000010000";
wait for Clk_period;
Addr <= "0001000101100";
Trees_din <= "00000010000000000001011000001000";
wait for Clk_period;
Addr <= "0001000101101";
Trees_din <= "00000100000000000001011100000100";
wait for Clk_period;
Addr <= "0001000101110";
Trees_din <= "00000000001011100000101000100001";
wait for Clk_period;
Addr <= "0001000101111";
Trees_din <= "00000000010000100000101000100001";
wait for Clk_period;
Addr <= "0001000110000";
Trees_din <= "00000101000000000000000000000100";
wait for Clk_period;
Addr <= "0001000110001";
Trees_din <= "00000000000110010000101000100001";
wait for Clk_period;
Addr <= "0001000110010";
Trees_din <= "00000000000101100000101000100001";
wait for Clk_period;
Addr <= "0001000110011";
Trees_din <= "00000010000000000001001000001000";
wait for Clk_period;
Addr <= "0001000110100";
Trees_din <= "00000110000000000101111000000100";
wait for Clk_period;
Addr <= "0001000110101";
Trees_din <= "00000000010111000000101000100001";
wait for Clk_period;
Addr <= "0001000110110";
Trees_din <= "00000000010100000000101000100001";
wait for Clk_period;
Addr <= "0001000110111";
Trees_din <= "00000010000000000100100100000100";
wait for Clk_period;
Addr <= "0001000111000";
Trees_din <= "00000000000111110000101000100001";
wait for Clk_period;
Addr <= "0001000111001";
Trees_din <= "00000000000001000000101000100001";
wait for Clk_period;
Addr <= "0001000111010";
Trees_din <= "00000111000000000010101000010000";
wait for Clk_period;
Addr <= "0001000111011";
Trees_din <= "00000001000000000000001000001000";
wait for Clk_period;
Addr <= "0001000111100";
Trees_din <= "00000001000000000101110000000100";
wait for Clk_period;
Addr <= "0001000111101";
Trees_din <= "00000000001110000000101000100001";
wait for Clk_period;
Addr <= "0001000111110";
Trees_din <= "00000000001101000000101000100001";
wait for Clk_period;
Addr <= "0001000111111";
Trees_din <= "00000101000000000101011100000100";
wait for Clk_period;
Addr <= "0001001000000";
Trees_din <= "00000000000100100000101000100001";
wait for Clk_period;
Addr <= "0001001000001";
Trees_din <= "00000000010111000000101000100001";
wait for Clk_period;
Addr <= "0001001000010";
Trees_din <= "00000110000000000000111100001000";
wait for Clk_period;
Addr <= "0001001000011";
Trees_din <= "00000010000000000000101000000100";
wait for Clk_period;
Addr <= "0001001000100";
Trees_din <= "00000000010000010000101000100001";
wait for Clk_period;
Addr <= "0001001000101";
Trees_din <= "00000000000110110000101000100001";
wait for Clk_period;
Addr <= "0001001000110";
Trees_din <= "00000111000000000101010000000100";
wait for Clk_period;
Addr <= "0001001000111";
Trees_din <= "00000000010000110000101000100001";
wait for Clk_period;
Addr <= "0001001001000";
Trees_din <= "00000000010100000000101000100001";
wait for Clk_period;
Addr <= "0001001001001";
Trees_din <= "00000111000000000010100101000000";
wait for Clk_period;
Addr <= "0001001001010";
Trees_din <= "00000010000000000101001000100000";
wait for Clk_period;
Addr <= "0001001001011";
Trees_din <= "00000100000000000101100000010000";
wait for Clk_period;
Addr <= "0001001001100";
Trees_din <= "00000111000000000000001000001000";
wait for Clk_period;
Addr <= "0001001001101";
Trees_din <= "00000110000000000011001100000100";
wait for Clk_period;
Addr <= "0001001001110";
Trees_din <= "00000000001111110000101000100001";
wait for Clk_period;
Addr <= "0001001001111";
Trees_din <= "00000000000000110000101000100001";
wait for Clk_period;
Addr <= "0001001010000";
Trees_din <= "00000000000000000000111100000100";
wait for Clk_period;
Addr <= "0001001010001";
Trees_din <= "00000000000001000000101000100001";
wait for Clk_period;
Addr <= "0001001010010";
Trees_din <= "00000000010110010000101000100001";
wait for Clk_period;
Addr <= "0001001010011";
Trees_din <= "00000011000000000010111100001000";
wait for Clk_period;
Addr <= "0001001010100";
Trees_din <= "00000011000000000101101100000100";
wait for Clk_period;
Addr <= "0001001010101";
Trees_din <= "00000000000100000000101000100001";
wait for Clk_period;
Addr <= "0001001010110";
Trees_din <= "00000000001001100000101000100001";
wait for Clk_period;
Addr <= "0001001010111";
Trees_din <= "00000100000000000110010000000100";
wait for Clk_period;
Addr <= "0001001011000";
Trees_din <= "00000000001010100000101000100001";
wait for Clk_period;
Addr <= "0001001011001";
Trees_din <= "00000000000110100000101000100001";
wait for Clk_period;
Addr <= "0001001011010";
Trees_din <= "00000100000000000011000000010000";
wait for Clk_period;
Addr <= "0001001011011";
Trees_din <= "00000101000000000001100000001000";
wait for Clk_period;
Addr <= "0001001011100";
Trees_din <= "00000010000000000100000100000100";
wait for Clk_period;
Addr <= "0001001011101";
Trees_din <= "00000000001101100000101000100001";
wait for Clk_period;
Addr <= "0001001011110";
Trees_din <= "00000000001111000000101000100001";
wait for Clk_period;
Addr <= "0001001011111";
Trees_din <= "00000000000000000100111000000100";
wait for Clk_period;
Addr <= "0001001100000";
Trees_din <= "00000000010101110000101000100001";
wait for Clk_period;
Addr <= "0001001100001";
Trees_din <= "00000000001011010000101000100001";
wait for Clk_period;
Addr <= "0001001100010";
Trees_din <= "00000000000000000011011000001000";
wait for Clk_period;
Addr <= "0001001100011";
Trees_din <= "00000111000000000000000000000100";
wait for Clk_period;
Addr <= "0001001100100";
Trees_din <= "00000000001111110000101000100001";
wait for Clk_period;
Addr <= "0001001100101";
Trees_din <= "00000000001001100000101000100001";
wait for Clk_period;
Addr <= "0001001100110";
Trees_din <= "00000000000000000000101000000100";
wait for Clk_period;
Addr <= "0001001100111";
Trees_din <= "00000000000000010000101000100001";
wait for Clk_period;
Addr <= "0001001101000";
Trees_din <= "00000000010010010000101000100001";
wait for Clk_period;
Addr <= "0001001101001";
Trees_din <= "00000111000000000100111100100000";
wait for Clk_period;
Addr <= "0001001101010";
Trees_din <= "00000001000000000011000000010000";
wait for Clk_period;
Addr <= "0001001101011";
Trees_din <= "00000110000000000000000000001000";
wait for Clk_period;
Addr <= "0001001101100";
Trees_din <= "00000011000000000010010100000100";
wait for Clk_period;
Addr <= "0001001101101";
Trees_din <= "00000000010110110000101000100001";
wait for Clk_period;
Addr <= "0001001101110";
Trees_din <= "00000000010110010000101000100001";
wait for Clk_period;
Addr <= "0001001101111";
Trees_din <= "00000100000000000000110100000100";
wait for Clk_period;
Addr <= "0001001110000";
Trees_din <= "00000000000011110000101000100001";
wait for Clk_period;
Addr <= "0001001110001";
Trees_din <= "00000000001010100000101000100001";
wait for Clk_period;
Addr <= "0001001110010";
Trees_din <= "00000001000000000010100000001000";
wait for Clk_period;
Addr <= "0001001110011";
Trees_din <= "00000110000000000100011100000100";
wait for Clk_period;
Addr <= "0001001110100";
Trees_din <= "00000000010011110000101000100001";
wait for Clk_period;
Addr <= "0001001110101";
Trees_din <= "00000000010100010000101000100001";
wait for Clk_period;
Addr <= "0001001110110";
Trees_din <= "00000100000000000000101100000100";
wait for Clk_period;
Addr <= "0001001110111";
Trees_din <= "00000000010100110000101000100001";
wait for Clk_period;
Addr <= "0001001111000";
Trees_din <= "00000000000111110000101000100001";
wait for Clk_period;
Addr <= "0001001111001";
Trees_din <= "00000111000000000100000000010000";
wait for Clk_period;
Addr <= "0001001111010";
Trees_din <= "00000010000000000101101000001000";
wait for Clk_period;
Addr <= "0001001111011";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "0001001111100";
Trees_din <= "00000000000111110000101000100001";
wait for Clk_period;
Addr <= "0001001111101";
Trees_din <= "00000000000101110000101000100001";
wait for Clk_period;
Addr <= "0001001111110";
Trees_din <= "00000101000000000101111100000100";
wait for Clk_period;
Addr <= "0001001111111";
Trees_din <= "00000000001010010000101000100001";
wait for Clk_period;
Addr <= "0001010000000";
Trees_din <= "00000000001010000000101000100001";
wait for Clk_period;
Addr <= "0001010000001";
Trees_din <= "00000110000000000010101100001000";
wait for Clk_period;
Addr <= "0001010000010";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "0001010000011";
Trees_din <= "00000000000111000000101000100001";
wait for Clk_period;
Addr <= "0001010000100";
Trees_din <= "00000000000001110000101000100001";
wait for Clk_period;
Addr <= "0001010000101";
Trees_din <= "00000110000000000001111100000100";
wait for Clk_period;
Addr <= "0001010000110";
Trees_din <= "00000000010111010000101000100001";
wait for Clk_period;
Addr <= "0001010000111";
Trees_din <= "00000000000100000000101000100001";
wait for Clk_period;



----------tree 5-------------------

Addr <= "0001010001000";
Trees_din <= "00000010000000000101011110000000";
wait for Clk_period;
Addr <= "0001010001001";
Trees_din <= "00000011000000000011111001000000";
wait for Clk_period;
Addr <= "0001010001010";
Trees_din <= "00000000000000000100110000100000";
wait for Clk_period;
Addr <= "0001010001011";
Trees_din <= "00000100000000000000000100010000";
wait for Clk_period;
Addr <= "0001010001100";
Trees_din <= "00000010000000000011110100001000";
wait for Clk_period;
Addr <= "0001010001101";
Trees_din <= "00000110000000000011110100000100";
wait for Clk_period;
Addr <= "0001010001110";
Trees_din <= "00000000011000110000000000000011";
wait for Clk_period;
Addr <= "0001010001111";
Trees_din <= "00000000001111100000000000000011";
wait for Clk_period;
Addr <= "0001010010000";
Trees_din <= "00000100000000000010000100000100";
wait for Clk_period;
Addr <= "0001010010001";
Trees_din <= "00000000001110010000000000000011";
wait for Clk_period;
Addr <= "0001010010010";
Trees_din <= "00000000000101010000000000000011";
wait for Clk_period;
Addr <= "0001010010011";
Trees_din <= "00000101000000000011110100001000";
wait for Clk_period;
Addr <= "0001010010100";
Trees_din <= "00000001000000000010101100000100";
wait for Clk_period;
Addr <= "0001010010101";
Trees_din <= "00000000000011000000000000000011";
wait for Clk_period;
Addr <= "0001010010110";
Trees_din <= "00000000010001110000000000000011";
wait for Clk_period;
Addr <= "0001010010111";
Trees_din <= "00000110000000000100001100000100";
wait for Clk_period;
Addr <= "0001010011000";
Trees_din <= "00000000001001000000000000000011";
wait for Clk_period;
Addr <= "0001010011001";
Trees_din <= "00000000001101010000000000000011";
wait for Clk_period;
Addr <= "0001010011010";
Trees_din <= "00000010000000000010010100010000";
wait for Clk_period;
Addr <= "0001010011011";
Trees_din <= "00000101000000000000110000001000";
wait for Clk_period;
Addr <= "0001010011100";
Trees_din <= "00000111000000000010111100000100";
wait for Clk_period;
Addr <= "0001010011101";
Trees_din <= "00000000001011110000000000000011";
wait for Clk_period;
Addr <= "0001010011110";
Trees_din <= "00000000000101100000000000000011";
wait for Clk_period;
Addr <= "0001010011111";
Trees_din <= "00000011000000000010100100000100";
wait for Clk_period;
Addr <= "0001010100000";
Trees_din <= "00000000010000010000000000000011";
wait for Clk_period;
Addr <= "0001010100001";
Trees_din <= "00000000000110000000000000000011";
wait for Clk_period;
Addr <= "0001010100010";
Trees_din <= "00000100000000000010001100001000";
wait for Clk_period;
Addr <= "0001010100011";
Trees_din <= "00000001000000000110000100000100";
wait for Clk_period;
Addr <= "0001010100100";
Trees_din <= "00000000001101000000000000000011";
wait for Clk_period;
Addr <= "0001010100101";
Trees_din <= "00000000010101100000000000000011";
wait for Clk_period;
Addr <= "0001010100110";
Trees_din <= "00000001000000000001101100000100";
wait for Clk_period;
Addr <= "0001010100111";
Trees_din <= "00000000001011100000000000000011";
wait for Clk_period;
Addr <= "0001010101000";
Trees_din <= "00000000001111010000000000000011";
wait for Clk_period;
Addr <= "0001010101001";
Trees_din <= "00000010000000000101000100100000";
wait for Clk_period;
Addr <= "0001010101010";
Trees_din <= "00000100000000000000110100010000";
wait for Clk_period;
Addr <= "0001010101011";
Trees_din <= "00000111000000000000011000001000";
wait for Clk_period;
Addr <= "0001010101100";
Trees_din <= "00000110000000000110010000000100";
wait for Clk_period;
Addr <= "0001010101101";
Trees_din <= "00000000010010110000000000000011";
wait for Clk_period;
Addr <= "0001010101110";
Trees_din <= "00000000001100000000000000000011";
wait for Clk_period;
Addr <= "0001010101111";
Trees_din <= "00000111000000000100111100000100";
wait for Clk_period;
Addr <= "0001010110000";
Trees_din <= "00000000001010000000000000000011";
wait for Clk_period;
Addr <= "0001010110001";
Trees_din <= "00000000001110000000000000000011";
wait for Clk_period;
Addr <= "0001010110010";
Trees_din <= "00000010000000000010011000001000";
wait for Clk_period;
Addr <= "0001010110011";
Trees_din <= "00000010000000000000100000000100";
wait for Clk_period;
Addr <= "0001010110100";
Trees_din <= "00000000001000110000000000000011";
wait for Clk_period;
Addr <= "0001010110101";
Trees_din <= "00000000010100010000000000000011";
wait for Clk_period;
Addr <= "0001010110110";
Trees_din <= "00000000000000000001001000000100";
wait for Clk_period;
Addr <= "0001010110111";
Trees_din <= "00000000010001000000000000000011";
wait for Clk_period;
Addr <= "0001010111000";
Trees_din <= "00000000010100100000000000000011";
wait for Clk_period;
Addr <= "0001010111001";
Trees_din <= "00000101000000000010001000010000";
wait for Clk_period;
Addr <= "0001010111010";
Trees_din <= "00000011000000000000010100001000";
wait for Clk_period;
Addr <= "0001010111011";
Trees_din <= "00000100000000000100100100000100";
wait for Clk_period;
Addr <= "0001010111100";
Trees_din <= "00000000001110110000000000000011";
wait for Clk_period;
Addr <= "0001010111101";
Trees_din <= "00000000000111000000000000000011";
wait for Clk_period;
Addr <= "0001010111110";
Trees_din <= "00000010000000000100111100000100";
wait for Clk_period;
Addr <= "0001010111111";
Trees_din <= "00000000001111010000000000000011";
wait for Clk_period;
Addr <= "0001011000000";
Trees_din <= "00000000000011100000000000000011";
wait for Clk_period;
Addr <= "0001011000001";
Trees_din <= "00000100000000000011101100001000";
wait for Clk_period;
Addr <= "0001011000010";
Trees_din <= "00000111000000000011011100000100";
wait for Clk_period;
Addr <= "0001011000011";
Trees_din <= "00000000010010100000000000000011";
wait for Clk_period;
Addr <= "0001011000100";
Trees_din <= "00000000000110000000000000000011";
wait for Clk_period;
Addr <= "0001011000101";
Trees_din <= "00000111000000000100111000000100";
wait for Clk_period;
Addr <= "0001011000110";
Trees_din <= "00000000001111100000000000000011";
wait for Clk_period;
Addr <= "0001011000111";
Trees_din <= "00000000010111000000000000000011";
wait for Clk_period;
Addr <= "0001011001000";
Trees_din <= "00000010000000000011100001000000";
wait for Clk_period;
Addr <= "0001011001001";
Trees_din <= "00000000000000000010111000100000";
wait for Clk_period;
Addr <= "0001011001010";
Trees_din <= "00000100000000000101110100010000";
wait for Clk_period;
Addr <= "0001011001011";
Trees_din <= "00000011000000000110010000001000";
wait for Clk_period;
Addr <= "0001011001100";
Trees_din <= "00000010000000000011001000000100";
wait for Clk_period;
Addr <= "0001011001101";
Trees_din <= "00000000001000100000000000000011";
wait for Clk_period;
Addr <= "0001011001110";
Trees_din <= "00000000010010100000000000000011";
wait for Clk_period;
Addr <= "0001011001111";
Trees_din <= "00000001000000000000000100000100";
wait for Clk_period;
Addr <= "0001011010000";
Trees_din <= "00000000010000100000000000000011";
wait for Clk_period;
Addr <= "0001011010001";
Trees_din <= "00000000000110010000000000000011";
wait for Clk_period;
Addr <= "0001011010010";
Trees_din <= "00000110000000000001000000001000";
wait for Clk_period;
Addr <= "0001011010011";
Trees_din <= "00000110000000000001001100000100";
wait for Clk_period;
Addr <= "0001011010100";
Trees_din <= "00000000010100100000000000000011";
wait for Clk_period;
Addr <= "0001011010101";
Trees_din <= "00000000010100010000000000000011";
wait for Clk_period;
Addr <= "0001011010110";
Trees_din <= "00000101000000000101010100000100";
wait for Clk_period;
Addr <= "0001011010111";
Trees_din <= "00000000001010000000000000000011";
wait for Clk_period;
Addr <= "0001011011000";
Trees_din <= "00000000001001100000000000000011";
wait for Clk_period;
Addr <= "0001011011001";
Trees_din <= "00000010000000000000110100010000";
wait for Clk_period;
Addr <= "0001011011010";
Trees_din <= "00000111000000000100101100001000";
wait for Clk_period;
Addr <= "0001011011011";
Trees_din <= "00000100000000000101110000000100";
wait for Clk_period;
Addr <= "0001011011100";
Trees_din <= "00000000001010000000000000000011";
wait for Clk_period;
Addr <= "0001011011101";
Trees_din <= "00000000000101100000000000000011";
wait for Clk_period;
Addr <= "0001011011110";
Trees_din <= "00000100000000000110010000000100";
wait for Clk_period;
Addr <= "0001011011111";
Trees_din <= "00000000000101000000000000000011";
wait for Clk_period;
Addr <= "0001011100000";
Trees_din <= "00000000001101100000000000000011";
wait for Clk_period;
Addr <= "0001011100001";
Trees_din <= "00000110000000000100101100001000";
wait for Clk_period;
Addr <= "0001011100010";
Trees_din <= "00000000000000000000000100000100";
wait for Clk_period;
Addr <= "0001011100011";
Trees_din <= "00000000000010110000000000000011";
wait for Clk_period;
Addr <= "0001011100100";
Trees_din <= "00000000000110110000000000000011";
wait for Clk_period;
Addr <= "0001011100101";
Trees_din <= "00000001000000000011110100000100";
wait for Clk_period;
Addr <= "0001011100110";
Trees_din <= "00000000000111000000000000000011";
wait for Clk_period;
Addr <= "0001011100111";
Trees_din <= "00000000000100100000000000000011";
wait for Clk_period;
Addr <= "0001011101000";
Trees_din <= "00000100000000000011000000100000";
wait for Clk_period;
Addr <= "0001011101001";
Trees_din <= "00000000000000000000100000010000";
wait for Clk_period;
Addr <= "0001011101010";
Trees_din <= "00000110000000000000100000001000";
wait for Clk_period;
Addr <= "0001011101011";
Trees_din <= "00000011000000000011000100000100";
wait for Clk_period;
Addr <= "0001011101100";
Trees_din <= "00000000000010000000000000000011";
wait for Clk_period;
Addr <= "0001011101101";
Trees_din <= "00000000010010110000000000000011";
wait for Clk_period;
Addr <= "0001011101110";
Trees_din <= "00000101000000000101011100000100";
wait for Clk_period;
Addr <= "0001011101111";
Trees_din <= "00000000000101010000000000000011";
wait for Clk_period;
Addr <= "0001011110000";
Trees_din <= "00000000001111010000000000000011";
wait for Clk_period;
Addr <= "0001011110001";
Trees_din <= "00000001000000000000111000001000";
wait for Clk_period;
Addr <= "0001011110010";
Trees_din <= "00000011000000000011101100000100";
wait for Clk_period;
Addr <= "0001011110011";
Trees_din <= "00000000010010110000000000000011";
wait for Clk_period;
Addr <= "0001011110100";
Trees_din <= "00000000010101000000000000000011";
wait for Clk_period;
Addr <= "0001011110101";
Trees_din <= "00000001000000000001000100000100";
wait for Clk_period;
Addr <= "0001011110110";
Trees_din <= "00000000000110010000000000000011";
wait for Clk_period;
Addr <= "0001011110111";
Trees_din <= "00000000001001100000000000000011";
wait for Clk_period;
Addr <= "0001011111000";
Trees_din <= "00000111000000000010100000010000";
wait for Clk_period;
Addr <= "0001011111001";
Trees_din <= "00000110000000000010110000001000";
wait for Clk_period;
Addr <= "0001011111010";
Trees_din <= "00000000000000000000110000000100";
wait for Clk_period;
Addr <= "0001011111011";
Trees_din <= "00000000001010010000000000000011";
wait for Clk_period;
Addr <= "0001011111100";
Trees_din <= "00000000001011100000000000000011";
wait for Clk_period;
Addr <= "0001011111101";
Trees_din <= "00000011000000000101111100000100";
wait for Clk_period;
Addr <= "0001011111110";
Trees_din <= "00000000000000010000000000000011";
wait for Clk_period;
Addr <= "0001011111111";
Trees_din <= "00000000010010110000000000000011";
wait for Clk_period;
Addr <= "0001100000000";
Trees_din <= "00000000000000000011010100001000";
wait for Clk_period;
Addr <= "0001100000001";
Trees_din <= "00000100000000000100111100000100";
wait for Clk_period;
Addr <= "0001100000010";
Trees_din <= "00000000000001100000000000000011";
wait for Clk_period;
Addr <= "0001100000011";
Trees_din <= "00000000001001000000000000000011";
wait for Clk_period;
Addr <= "0001100000100";
Trees_din <= "00000111000000000110000000000100";
wait for Clk_period;
Addr <= "0001100000101";
Trees_din <= "00000000001101100000000000000011";
wait for Clk_period;
Addr <= "0001100000110";
Trees_din <= "00000000011000110000000000000011";
wait for Clk_period;



----------tree 6-------------------

Addr <= "0001100000111";
Trees_din <= "00000010000000000010111010000000";
wait for Clk_period;
Addr <= "0001100001000";
Trees_din <= "00000010000000000001001101000000";
wait for Clk_period;
Addr <= "0001100001001";
Trees_din <= "00000010000000000011011100100000";
wait for Clk_period;
Addr <= "0001100001010";
Trees_din <= "00000001000000000100011100010000";
wait for Clk_period;
Addr <= "0001100001011";
Trees_din <= "00000011000000000010001000001000";
wait for Clk_period;
Addr <= "0001100001100";
Trees_din <= "00000010000000000100000000000100";
wait for Clk_period;
Addr <= "0001100001101";
Trees_din <= "00000000001011110000111000011001";
wait for Clk_period;
Addr <= "0001100001110";
Trees_din <= "00000000001011000000111000011001";
wait for Clk_period;
Addr <= "0001100001111";
Trees_din <= "00000101000000000011001100000100";
wait for Clk_period;
Addr <= "0001100010000";
Trees_din <= "00000000001100000000111000011001";
wait for Clk_period;
Addr <= "0001100010001";
Trees_din <= "00000000000111000000111000011001";
wait for Clk_period;
Addr <= "0001100010010";
Trees_din <= "00000101000000000110001000001000";
wait for Clk_period;
Addr <= "0001100010011";
Trees_din <= "00000100000000000000000000000100";
wait for Clk_period;
Addr <= "0001100010100";
Trees_din <= "00000000001000100000111000011001";
wait for Clk_period;
Addr <= "0001100010101";
Trees_din <= "00000000000000100000111000011001";
wait for Clk_period;
Addr <= "0001100010110";
Trees_din <= "00000001000000000001001000000100";
wait for Clk_period;
Addr <= "0001100010111";
Trees_din <= "00000000001000000000111000011001";
wait for Clk_period;
Addr <= "0001100011000";
Trees_din <= "00000000000111100000111000011001";
wait for Clk_period;
Addr <= "0001100011001";
Trees_din <= "00000111000000000010001000010000";
wait for Clk_period;
Addr <= "0001100011010";
Trees_din <= "00000100000000000011010000001000";
wait for Clk_period;
Addr <= "0001100011011";
Trees_din <= "00000100000000000000000100000100";
wait for Clk_period;
Addr <= "0001100011100";
Trees_din <= "00000000001000110000111000011001";
wait for Clk_period;
Addr <= "0001100011101";
Trees_din <= "00000000010000000000111000011001";
wait for Clk_period;
Addr <= "0001100011110";
Trees_din <= "00000011000000000100010100000100";
wait for Clk_period;
Addr <= "0001100011111";
Trees_din <= "00000000000111100000111000011001";
wait for Clk_period;
Addr <= "0001100100000";
Trees_din <= "00000000011000000000111000011001";
wait for Clk_period;
Addr <= "0001100100001";
Trees_din <= "00000100000000000010111000001000";
wait for Clk_period;
Addr <= "0001100100010";
Trees_din <= "00000100000000000010000100000100";
wait for Clk_period;
Addr <= "0001100100011";
Trees_din <= "00000000000010110000111000011001";
wait for Clk_period;
Addr <= "0001100100100";
Trees_din <= "00000000000000100000111000011001";
wait for Clk_period;
Addr <= "0001100100101";
Trees_din <= "00000111000000000001001000000100";
wait for Clk_period;
Addr <= "0001100100110";
Trees_din <= "00000000010010110000111000011001";
wait for Clk_period;
Addr <= "0001100100111";
Trees_din <= "00000000001101110000111000011001";
wait for Clk_period;
Addr <= "0001100101000";
Trees_din <= "00000110000000000101111000100000";
wait for Clk_period;
Addr <= "0001100101001";
Trees_din <= "00000010000000000100010100010000";
wait for Clk_period;
Addr <= "0001100101010";
Trees_din <= "00000010000000000101000000001000";
wait for Clk_period;
Addr <= "0001100101011";
Trees_din <= "00000001000000000110000000000100";
wait for Clk_period;
Addr <= "0001100101100";
Trees_din <= "00000000001101100000111000011001";
wait for Clk_period;
Addr <= "0001100101101";
Trees_din <= "00000000010100010000111000011001";
wait for Clk_period;
Addr <= "0001100101110";
Trees_din <= "00000111000000000100101100000100";
wait for Clk_period;
Addr <= "0001100101111";
Trees_din <= "00000000001100000000111000011001";
wait for Clk_period;
Addr <= "0001100110000";
Trees_din <= "00000000010101010000111000011001";
wait for Clk_period;
Addr <= "0001100110001";
Trees_din <= "00000111000000000001110000001000";
wait for Clk_period;
Addr <= "0001100110010";
Trees_din <= "00000100000000000101110100000100";
wait for Clk_period;
Addr <= "0001100110011";
Trees_din <= "00000000000111000000111000011001";
wait for Clk_period;
Addr <= "0001100110100";
Trees_din <= "00000000000110110000111000011001";
wait for Clk_period;
Addr <= "0001100110101";
Trees_din <= "00000010000000000100011100000100";
wait for Clk_period;
Addr <= "0001100110110";
Trees_din <= "00000000000111000000111000011001";
wait for Clk_period;
Addr <= "0001100110111";
Trees_din <= "00000000001101000000111000011001";
wait for Clk_period;
Addr <= "0001100111000";
Trees_din <= "00000100000000000100100100010000";
wait for Clk_period;
Addr <= "0001100111001";
Trees_din <= "00000011000000000001011000001000";
wait for Clk_period;
Addr <= "0001100111010";
Trees_din <= "00000001000000000000000000000100";
wait for Clk_period;
Addr <= "0001100111011";
Trees_din <= "00000000001011000000111000011001";
wait for Clk_period;
Addr <= "0001100111100";
Trees_din <= "00000000010110000000111000011001";
wait for Clk_period;
Addr <= "0001100111101";
Trees_din <= "00000110000000000100010100000100";
wait for Clk_period;
Addr <= "0001100111110";
Trees_din <= "00000000000101000000111000011001";
wait for Clk_period;
Addr <= "0001100111111";
Trees_din <= "00000000000110000000111000011001";
wait for Clk_period;
Addr <= "0001101000000";
Trees_din <= "00000101000000000100101100001000";
wait for Clk_period;
Addr <= "0001101000001";
Trees_din <= "00000101000000000000110000000100";
wait for Clk_period;
Addr <= "0001101000010";
Trees_din <= "00000000010001100000111000011001";
wait for Clk_period;
Addr <= "0001101000011";
Trees_din <= "00000000000110100000111000011001";
wait for Clk_period;
Addr <= "0001101000100";
Trees_din <= "00000101000000000101001100000100";
wait for Clk_period;
Addr <= "0001101000101";
Trees_din <= "00000000011000110000111000011001";
wait for Clk_period;
Addr <= "0001101000110";
Trees_din <= "00000000000111010000111000011001";
wait for Clk_period;
Addr <= "0001101000111";
Trees_din <= "00000011000000000000111001000000";
wait for Clk_period;
Addr <= "0001101001000";
Trees_din <= "00000000000000000101111100100000";
wait for Clk_period;
Addr <= "0001101001001";
Trees_din <= "00000100000000000001011000010000";
wait for Clk_period;
Addr <= "0001101001010";
Trees_din <= "00000100000000000010010100001000";
wait for Clk_period;
Addr <= "0001101001011";
Trees_din <= "00000000000000000100001100000100";
wait for Clk_period;
Addr <= "0001101001100";
Trees_din <= "00000000000101000000111000011001";
wait for Clk_period;
Addr <= "0001101001101";
Trees_din <= "00000000001000110000111000011001";
wait for Clk_period;
Addr <= "0001101001110";
Trees_din <= "00000110000000000000110100000100";
wait for Clk_period;
Addr <= "0001101001111";
Trees_din <= "00000000000001110000111000011001";
wait for Clk_period;
Addr <= "0001101010000";
Trees_din <= "00000000010110110000111000011001";
wait for Clk_period;
Addr <= "0001101010001";
Trees_din <= "00000010000000000011010000001000";
wait for Clk_period;
Addr <= "0001101010010";
Trees_din <= "00000111000000000101111100000100";
wait for Clk_period;
Addr <= "0001101010011";
Trees_din <= "00000000010111100000111000011001";
wait for Clk_period;
Addr <= "0001101010100";
Trees_din <= "00000000001110010000111000011001";
wait for Clk_period;
Addr <= "0001101010101";
Trees_din <= "00000100000000000110000000000100";
wait for Clk_period;
Addr <= "0001101010110";
Trees_din <= "00000000000110100000111000011001";
wait for Clk_period;
Addr <= "0001101010111";
Trees_din <= "00000000000010010000111000011001";
wait for Clk_period;
Addr <= "0001101011000";
Trees_din <= "00000000000000000001100000010000";
wait for Clk_period;
Addr <= "0001101011001";
Trees_din <= "00000101000000000100000100001000";
wait for Clk_period;
Addr <= "0001101011010";
Trees_din <= "00000011000000000000000100000100";
wait for Clk_period;
Addr <= "0001101011011";
Trees_din <= "00000000000000000000111000011001";
wait for Clk_period;
Addr <= "0001101011100";
Trees_din <= "00000000011000000000111000011001";
wait for Clk_period;
Addr <= "0001101011101";
Trees_din <= "00000010000000000100001000000100";
wait for Clk_period;
Addr <= "0001101011110";
Trees_din <= "00000000001100110000111000011001";
wait for Clk_period;
Addr <= "0001101011111";
Trees_din <= "00000000001101010000111000011001";
wait for Clk_period;
Addr <= "0001101100000";
Trees_din <= "00000001000000000011010100001000";
wait for Clk_period;
Addr <= "0001101100001";
Trees_din <= "00000101000000000100001000000100";
wait for Clk_period;
Addr <= "0001101100010";
Trees_din <= "00000000000000000000111000011001";
wait for Clk_period;
Addr <= "0001101100011";
Trees_din <= "00000000001111000000111000011001";
wait for Clk_period;
Addr <= "0001101100100";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "0001101100101";
Trees_din <= "00000000010010110000111000011001";
wait for Clk_period;
Addr <= "0001101100110";
Trees_din <= "00000000010100110000111000011001";
wait for Clk_period;
Addr <= "0001101100111";
Trees_din <= "00000110000000000000011000100000";
wait for Clk_period;
Addr <= "0001101101000";
Trees_din <= "00000100000000000011000100010000";
wait for Clk_period;
Addr <= "0001101101001";
Trees_din <= "00000100000000000001010100001000";
wait for Clk_period;
Addr <= "0001101101010";
Trees_din <= "00000111000000000000000000000100";
wait for Clk_period;
Addr <= "0001101101011";
Trees_din <= "00000000010111100000111000011001";
wait for Clk_period;
Addr <= "0001101101100";
Trees_din <= "00000000000010010000111000011001";
wait for Clk_period;
Addr <= "0001101101101";
Trees_din <= "00000101000000000011000000000100";
wait for Clk_period;
Addr <= "0001101101110";
Trees_din <= "00000000001011000000111000011001";
wait for Clk_period;
Addr <= "0001101101111";
Trees_din <= "00000000000110000000111000011001";
wait for Clk_period;
Addr <= "0001101110000";
Trees_din <= "00000100000000000001010100001000";
wait for Clk_period;
Addr <= "0001101110001";
Trees_din <= "00000010000000000001111000000100";
wait for Clk_period;
Addr <= "0001101110010";
Trees_din <= "00000000010101100000111000011001";
wait for Clk_period;
Addr <= "0001101110011";
Trees_din <= "00000000000001000000111000011001";
wait for Clk_period;
Addr <= "0001101110100";
Trees_din <= "00000101000000000100000100000100";
wait for Clk_period;
Addr <= "0001101110101";
Trees_din <= "00000000010111000000111000011001";
wait for Clk_period;
Addr <= "0001101110110";
Trees_din <= "00000000010001000000111000011001";
wait for Clk_period;
Addr <= "0001101110111";
Trees_din <= "00000011000000000101000000010000";
wait for Clk_period;
Addr <= "0001101111000";
Trees_din <= "00000100000000000010001000001000";
wait for Clk_period;
Addr <= "0001101111001";
Trees_din <= "00000101000000000101110000000100";
wait for Clk_period;
Addr <= "0001101111010";
Trees_din <= "00000000010111100000111000011001";
wait for Clk_period;
Addr <= "0001101111011";
Trees_din <= "00000000010111110000111000011001";
wait for Clk_period;
Addr <= "0001101111100";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "0001101111101";
Trees_din <= "00000000001111100000111000011001";
wait for Clk_period;
Addr <= "0001101111110";
Trees_din <= "00000000000111010000111000011001";
wait for Clk_period;
Addr <= "0001101111111";
Trees_din <= "00000011000000000000001100001000";
wait for Clk_period;
Addr <= "0001110000000";
Trees_din <= "00000101000000000101011100000100";
wait for Clk_period;
Addr <= "0001110000001";
Trees_din <= "00000000001011110000111000011001";
wait for Clk_period;
Addr <= "0001110000010";
Trees_din <= "00000000010000100000111000011001";
wait for Clk_period;
Addr <= "0001110000011";
Trees_din <= "00000001000000000001011000000100";
wait for Clk_period;
Addr <= "0001110000100";
Trees_din <= "00000000001010000000111000011001";
wait for Clk_period;
Addr <= "0001110000101";
Trees_din <= "00000000000101110000111000011001";
wait for Clk_period;



----------tree 7-------------------

Addr <= "0001110000110";
Trees_din <= "00000010000000000010111010000000";
wait for Clk_period;
Addr <= "0001110000111";
Trees_din <= "00000100000000000011110001000000";
wait for Clk_period;
Addr <= "0001110001000";
Trees_din <= "00000110000000000000011000100000";
wait for Clk_period;
Addr <= "0001110001001";
Trees_din <= "00000110000000000000010000010000";
wait for Clk_period;
Addr <= "0001110001010";
Trees_din <= "00000110000000000000110000001000";
wait for Clk_period;
Addr <= "0001110001011";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "0001110001100";
Trees_din <= "00000000001001000001000000010111";
wait for Clk_period;
Addr <= "0001110001101";
Trees_din <= "00000000000100000001000000010111";
wait for Clk_period;
Addr <= "0001110001110";
Trees_din <= "00000100000000000101100000000100";
wait for Clk_period;
Addr <= "0001110001111";
Trees_din <= "00000000000110010001000000010111";
wait for Clk_period;
Addr <= "0001110010000";
Trees_din <= "00000000001110100001000000010111";
wait for Clk_period;
Addr <= "0001110010001";
Trees_din <= "00000000000000000010001000001000";
wait for Clk_period;
Addr <= "0001110010010";
Trees_din <= "00000001000000000001100000000100";
wait for Clk_period;
Addr <= "0001110010011";
Trees_din <= "00000000000011110001000000010111";
wait for Clk_period;
Addr <= "0001110010100";
Trees_din <= "00000000010100100001000000010111";
wait for Clk_period;
Addr <= "0001110010101";
Trees_din <= "00000000000000000110001100000100";
wait for Clk_period;
Addr <= "0001110010110";
Trees_din <= "00000000000001110001000000010111";
wait for Clk_period;
Addr <= "0001110010111";
Trees_din <= "00000000010001000001000000010111";
wait for Clk_period;
Addr <= "0001110011000";
Trees_din <= "00000000000000000011010100010000";
wait for Clk_period;
Addr <= "0001110011001";
Trees_din <= "00000110000000000001100000001000";
wait for Clk_period;
Addr <= "0001110011010";
Trees_din <= "00000011000000000100000000000100";
wait for Clk_period;
Addr <= "0001110011011";
Trees_din <= "00000000010010010001000000010111";
wait for Clk_period;
Addr <= "0001110011100";
Trees_din <= "00000000000000100001000000010111";
wait for Clk_period;
Addr <= "0001110011101";
Trees_din <= "00000111000000000001001000000100";
wait for Clk_period;
Addr <= "0001110011110";
Trees_din <= "00000000000000100001000000010111";
wait for Clk_period;
Addr <= "0001110011111";
Trees_din <= "00000000000001010001000000010111";
wait for Clk_period;
Addr <= "0001110100000";
Trees_din <= "00000110000000000101001000001000";
wait for Clk_period;
Addr <= "0001110100001";
Trees_din <= "00000001000000000010110000000100";
wait for Clk_period;
Addr <= "0001110100010";
Trees_din <= "00000000010000100001000000010111";
wait for Clk_period;
Addr <= "0001110100011";
Trees_din <= "00000000010000110001000000010111";
wait for Clk_period;
Addr <= "0001110100100";
Trees_din <= "00000111000000000100011100000100";
wait for Clk_period;
Addr <= "0001110100101";
Trees_din <= "00000000000000100001000000010111";
wait for Clk_period;
Addr <= "0001110100110";
Trees_din <= "00000000010100010001000000010111";
wait for Clk_period;
Addr <= "0001110100111";
Trees_din <= "00000000000000000100100100100000";
wait for Clk_period;
Addr <= "0001110101000";
Trees_din <= "00000011000000000000110100010000";
wait for Clk_period;
Addr <= "0001110101001";
Trees_din <= "00000010000000000011000000001000";
wait for Clk_period;
Addr <= "0001110101010";
Trees_din <= "00000000000000000110000000000100";
wait for Clk_period;
Addr <= "0001110101011";
Trees_din <= "00000000010011100001000000010111";
wait for Clk_period;
Addr <= "0001110101100";
Trees_din <= "00000000000010110001000000010111";
wait for Clk_period;
Addr <= "0001110101101";
Trees_din <= "00000010000000000010000100000100";
wait for Clk_period;
Addr <= "0001110101110";
Trees_din <= "00000000010111010001000000010111";
wait for Clk_period;
Addr <= "0001110101111";
Trees_din <= "00000000001111110001000000010111";
wait for Clk_period;
Addr <= "0001110110000";
Trees_din <= "00000010000000000000010100001000";
wait for Clk_period;
Addr <= "0001110110001";
Trees_din <= "00000100000000000010001100000100";
wait for Clk_period;
Addr <= "0001110110010";
Trees_din <= "00000000000100000001000000010111";
wait for Clk_period;
Addr <= "0001110110011";
Trees_din <= "00000000010000110001000000010111";
wait for Clk_period;
Addr <= "0001110110100";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "0001110110101";
Trees_din <= "00000000001101110001000000010111";
wait for Clk_period;
Addr <= "0001110110110";
Trees_din <= "00000000010101000001000000010111";
wait for Clk_period;
Addr <= "0001110110111";
Trees_din <= "00000010000000000001110000010000";
wait for Clk_period;
Addr <= "0001110111000";
Trees_din <= "00000101000000000110001000001000";
wait for Clk_period;
Addr <= "0001110111001";
Trees_din <= "00000001000000000000101100000100";
wait for Clk_period;
Addr <= "0001110111010";
Trees_din <= "00000000000001010001000000010111";
wait for Clk_period;
Addr <= "0001110111011";
Trees_din <= "00000000010001110001000000010111";
wait for Clk_period;
Addr <= "0001110111100";
Trees_din <= "00000111000000000100000100000100";
wait for Clk_period;
Addr <= "0001110111101";
Trees_din <= "00000000001011010001000000010111";
wait for Clk_period;
Addr <= "0001110111110";
Trees_din <= "00000000010110100001000000010111";
wait for Clk_period;
Addr <= "0001110111111";
Trees_din <= "00000000000000000010011000001000";
wait for Clk_period;
Addr <= "0001111000000";
Trees_din <= "00000010000000000100111100000100";
wait for Clk_period;
Addr <= "0001111000001";
Trees_din <= "00000000000000010001000000010111";
wait for Clk_period;
Addr <= "0001111000010";
Trees_din <= "00000000001111110001000000010111";
wait for Clk_period;
Addr <= "0001111000011";
Trees_din <= "00000001000000000110001100000100";
wait for Clk_period;
Addr <= "0001111000100";
Trees_din <= "00000000001101110001000000010111";
wait for Clk_period;
Addr <= "0001111000101";
Trees_din <= "00000000000010010001000000010111";
wait for Clk_period;
Addr <= "0001111000110";
Trees_din <= "00000110000000000010100101000000";
wait for Clk_period;
Addr <= "0001111000111";
Trees_din <= "00000110000000000100110000100000";
wait for Clk_period;
Addr <= "0001111001000";
Trees_din <= "00000110000000000110000100010000";
wait for Clk_period;
Addr <= "0001111001001";
Trees_din <= "00000101000000000001011100001000";
wait for Clk_period;
Addr <= "0001111001010";
Trees_din <= "00000000000000000010001100000100";
wait for Clk_period;
Addr <= "0001111001011";
Trees_din <= "00000000010011110001000000010111";
wait for Clk_period;
Addr <= "0001111001100";
Trees_din <= "00000000000000100001000000010111";
wait for Clk_period;
Addr <= "0001111001101";
Trees_din <= "00000001000000000011101100000100";
wait for Clk_period;
Addr <= "0001111001110";
Trees_din <= "00000000001010110001000000010111";
wait for Clk_period;
Addr <= "0001111001111";
Trees_din <= "00000000001111110001000000010111";
wait for Clk_period;
Addr <= "0001111010000";
Trees_din <= "00000001000000000010010100001000";
wait for Clk_period;
Addr <= "0001111010001";
Trees_din <= "00000111000000000101110000000100";
wait for Clk_period;
Addr <= "0001111010010";
Trees_din <= "00000000001111100001000000010111";
wait for Clk_period;
Addr <= "0001111010011";
Trees_din <= "00000000011000110001000000010111";
wait for Clk_period;
Addr <= "0001111010100";
Trees_din <= "00000101000000000000100100000100";
wait for Clk_period;
Addr <= "0001111010101";
Trees_din <= "00000000010111110001000000010111";
wait for Clk_period;
Addr <= "0001111010110";
Trees_din <= "00000000010110000001000000010111";
wait for Clk_period;
Addr <= "0001111010111";
Trees_din <= "00000000000000000101000000010000";
wait for Clk_period;
Addr <= "0001111011000";
Trees_din <= "00000100000000000001100000001000";
wait for Clk_period;
Addr <= "0001111011001";
Trees_din <= "00000011000000000001000100000100";
wait for Clk_period;
Addr <= "0001111011010";
Trees_din <= "00000000000110000001000000010111";
wait for Clk_period;
Addr <= "0001111011011";
Trees_din <= "00000000010101000001000000010111";
wait for Clk_period;
Addr <= "0001111011100";
Trees_din <= "00000010000000000011100000000100";
wait for Clk_period;
Addr <= "0001111011101";
Trees_din <= "00000000010000000001000000010111";
wait for Clk_period;
Addr <= "0001111011110";
Trees_din <= "00000000001010010001000000010111";
wait for Clk_period;
Addr <= "0001111011111";
Trees_din <= "00000010000000000010001100001000";
wait for Clk_period;
Addr <= "0001111100000";
Trees_din <= "00000001000000000100110000000100";
wait for Clk_period;
Addr <= "0001111100001";
Trees_din <= "00000000001111010001000000010111";
wait for Clk_period;
Addr <= "0001111100010";
Trees_din <= "00000000010000100001000000010111";
wait for Clk_period;
Addr <= "0001111100011";
Trees_din <= "00000100000000000010110100000100";
wait for Clk_period;
Addr <= "0001111100100";
Trees_din <= "00000000010001010001000000010111";
wait for Clk_period;
Addr <= "0001111100101";
Trees_din <= "00000000001001010001000000010111";
wait for Clk_period;
Addr <= "0001111100110";
Trees_din <= "00000101000000000100110000100000";
wait for Clk_period;
Addr <= "0001111100111";
Trees_din <= "00000010000000000011100000010000";
wait for Clk_period;
Addr <= "0001111101000";
Trees_din <= "00000110000000000000001100001000";
wait for Clk_period;
Addr <= "0001111101001";
Trees_din <= "00000000000000000000001100000100";
wait for Clk_period;
Addr <= "0001111101010";
Trees_din <= "00000000001011000001000000010111";
wait for Clk_period;
Addr <= "0001111101011";
Trees_din <= "00000000000101110001000000010111";
wait for Clk_period;
Addr <= "0001111101100";
Trees_din <= "00000000000000000000100000000100";
wait for Clk_period;
Addr <= "0001111101101";
Trees_din <= "00000000000110000001000000010111";
wait for Clk_period;
Addr <= "0001111101110";
Trees_din <= "00000000010101100001000000010111";
wait for Clk_period;
Addr <= "0001111101111";
Trees_din <= "00000001000000000110010000001000";
wait for Clk_period;
Addr <= "0001111110000";
Trees_din <= "00000111000000000011101000000100";
wait for Clk_period;
Addr <= "0001111110001";
Trees_din <= "00000000001101000001000000010111";
wait for Clk_period;
Addr <= "0001111110010";
Trees_din <= "00000000000111000001000000010111";
wait for Clk_period;
Addr <= "0001111110011";
Trees_din <= "00000101000000000101101100000100";
wait for Clk_period;
Addr <= "0001111110100";
Trees_din <= "00000000000111000001000000010111";
wait for Clk_period;
Addr <= "0001111110101";
Trees_din <= "00000000001101000001000000010111";
wait for Clk_period;
Addr <= "0001111110110";
Trees_din <= "00000000000000000001111000010000";
wait for Clk_period;
Addr <= "0001111110111";
Trees_din <= "00000101000000000100100100001000";
wait for Clk_period;
Addr <= "0001111111000";
Trees_din <= "00000101000000000000111100000100";
wait for Clk_period;
Addr <= "0001111111001";
Trees_din <= "00000000010000110001000000010111";
wait for Clk_period;
Addr <= "0001111111010";
Trees_din <= "00000000000101000001000000010111";
wait for Clk_period;
Addr <= "0001111111011";
Trees_din <= "00000001000000000000110100000100";
wait for Clk_period;
Addr <= "0001111111100";
Trees_din <= "00000000001001000001000000010111";
wait for Clk_period;
Addr <= "0001111111101";
Trees_din <= "00000000010101100001000000010111";
wait for Clk_period;
Addr <= "0001111111110";
Trees_din <= "00000111000000000010011000001000";
wait for Clk_period;
Addr <= "0001111111111";
Trees_din <= "00000100000000000010000000000100";
wait for Clk_period;
Addr <= "0010000000000";
Trees_din <= "00000000010111000001000000010111";
wait for Clk_period;
Addr <= "0010000000001";
Trees_din <= "00000000000111000001000000010111";
wait for Clk_period;
Addr <= "0010000000010";
Trees_din <= "00000000000000000101001100000100";
wait for Clk_period;
Addr <= "0010000000011";
Trees_din <= "00000000000000100001000000010111";
wait for Clk_period;
Addr <= "0010000000100";
Trees_din <= "00000000001001110001000000010111";
wait for Clk_period;



----------tree 8-------------------

Addr <= "0010000000101";
Trees_din <= "00000010000000000011010010000000";
wait for Clk_period;
Addr <= "0010000000110";
Trees_din <= "00000101000000000011110001000000";
wait for Clk_period;
Addr <= "0010000000111";
Trees_din <= "00000000000000000011001100100000";
wait for Clk_period;
Addr <= "0010000001000";
Trees_din <= "00000110000000000000110100010000";
wait for Clk_period;
Addr <= "0010000001001";
Trees_din <= "00000011000000000011100000001000";
wait for Clk_period;
Addr <= "0010000001010";
Trees_din <= "00000011000000000010011100000100";
wait for Clk_period;
Addr <= "0010000001011";
Trees_din <= "00000000001110000001001000010001";
wait for Clk_period;
Addr <= "0010000001100";
Trees_din <= "00000000010001010001001000010001";
wait for Clk_period;
Addr <= "0010000001101";
Trees_din <= "00000001000000000010010100000100";
wait for Clk_period;
Addr <= "0010000001110";
Trees_din <= "00000000010100000001001000010001";
wait for Clk_period;
Addr <= "0010000001111";
Trees_din <= "00000000001011110001001000010001";
wait for Clk_period;
Addr <= "0010000010000";
Trees_din <= "00000110000000000101001100001000";
wait for Clk_period;
Addr <= "0010000010001";
Trees_din <= "00000101000000000010000100000100";
wait for Clk_period;
Addr <= "0010000010010";
Trees_din <= "00000000000001000001001000010001";
wait for Clk_period;
Addr <= "0010000010011";
Trees_din <= "00000000011000100001001000010001";
wait for Clk_period;
Addr <= "0010000010100";
Trees_din <= "00000101000000000001000100000100";
wait for Clk_period;
Addr <= "0010000010101";
Trees_din <= "00000000001110010001001000010001";
wait for Clk_period;
Addr <= "0010000010110";
Trees_din <= "00000000000111110001001000010001";
wait for Clk_period;
Addr <= "0010000010111";
Trees_din <= "00000011000000000100010100010000";
wait for Clk_period;
Addr <= "0010000011000";
Trees_din <= "00000100000000000100101100001000";
wait for Clk_period;
Addr <= "0010000011001";
Trees_din <= "00000100000000000101000000000100";
wait for Clk_period;
Addr <= "0010000011010";
Trees_din <= "00000000010101010001001000010001";
wait for Clk_period;
Addr <= "0010000011011";
Trees_din <= "00000000001001100001001000010001";
wait for Clk_period;
Addr <= "0010000011100";
Trees_din <= "00000100000000000000011100000100";
wait for Clk_period;
Addr <= "0010000011101";
Trees_din <= "00000000010101100001001000010001";
wait for Clk_period;
Addr <= "0010000011110";
Trees_din <= "00000000000111110001001000010001";
wait for Clk_period;
Addr <= "0010000011111";
Trees_din <= "00000010000000000011000000001000";
wait for Clk_period;
Addr <= "0010000100000";
Trees_din <= "00000010000000000101101000000100";
wait for Clk_period;
Addr <= "0010000100001";
Trees_din <= "00000000010000100001001000010001";
wait for Clk_period;
Addr <= "0010000100010";
Trees_din <= "00000000011000100001001000010001";
wait for Clk_period;
Addr <= "0010000100011";
Trees_din <= "00000110000000000010000100000100";
wait for Clk_period;
Addr <= "0010000100100";
Trees_din <= "00000000010101100001001000010001";
wait for Clk_period;
Addr <= "0010000100101";
Trees_din <= "00000000000110100001001000010001";
wait for Clk_period;
Addr <= "0010000100110";
Trees_din <= "00000010000000000001100000100000";
wait for Clk_period;
Addr <= "0010000100111";
Trees_din <= "00000010000000000000000000010000";
wait for Clk_period;
Addr <= "0010000101000";
Trees_din <= "00000010000000000010011100001000";
wait for Clk_period;
Addr <= "0010000101001";
Trees_din <= "00000110000000000001001100000100";
wait for Clk_period;
Addr <= "0010000101010";
Trees_din <= "00000000010111010001001000010001";
wait for Clk_period;
Addr <= "0010000101011";
Trees_din <= "00000000000110000001001000010001";
wait for Clk_period;
Addr <= "0010000101100";
Trees_din <= "00000100000000000010011000000100";
wait for Clk_period;
Addr <= "0010000101101";
Trees_din <= "00000000001100000001001000010001";
wait for Clk_period;
Addr <= "0010000101110";
Trees_din <= "00000000000111010001001000010001";
wait for Clk_period;
Addr <= "0010000101111";
Trees_din <= "00000101000000000001010000001000";
wait for Clk_period;
Addr <= "0010000110000";
Trees_din <= "00000001000000000010100100000100";
wait for Clk_period;
Addr <= "0010000110001";
Trees_din <= "00000000001010100001001000010001";
wait for Clk_period;
Addr <= "0010000110010";
Trees_din <= "00000000010010010001001000010001";
wait for Clk_period;
Addr <= "0010000110011";
Trees_din <= "00000111000000000010001100000100";
wait for Clk_period;
Addr <= "0010000110100";
Trees_din <= "00000000001101010001001000010001";
wait for Clk_period;
Addr <= "0010000110101";
Trees_din <= "00000000010001000001001000010001";
wait for Clk_period;
Addr <= "0010000110110";
Trees_din <= "00000001000000000101110100010000";
wait for Clk_period;
Addr <= "0010000110111";
Trees_din <= "00000010000000000001110100001000";
wait for Clk_period;
Addr <= "0010000111000";
Trees_din <= "00000100000000000001010000000100";
wait for Clk_period;
Addr <= "0010000111001";
Trees_din <= "00000000010001100001001000010001";
wait for Clk_period;
Addr <= "0010000111010";
Trees_din <= "00000000010001000001001000010001";
wait for Clk_period;
Addr <= "0010000111011";
Trees_din <= "00000010000000000010001100000100";
wait for Clk_period;
Addr <= "0010000111100";
Trees_din <= "00000000010001000001001000010001";
wait for Clk_period;
Addr <= "0010000111101";
Trees_din <= "00000000000011110001001000010001";
wait for Clk_period;
Addr <= "0010000111110";
Trees_din <= "00000100000000000001000100001000";
wait for Clk_period;
Addr <= "0010000111111";
Trees_din <= "00000010000000000100001100000100";
wait for Clk_period;
Addr <= "0010001000000";
Trees_din <= "00000000000000010001001000010001";
wait for Clk_period;
Addr <= "0010001000001";
Trees_din <= "00000000010111010001001000010001";
wait for Clk_period;
Addr <= "0010001000010";
Trees_din <= "00000100000000000100011100000100";
wait for Clk_period;
Addr <= "0010001000011";
Trees_din <= "00000000011000110001001000010001";
wait for Clk_period;
Addr <= "0010001000100";
Trees_din <= "00000000001010110001001000010001";
wait for Clk_period;
Addr <= "0010001000101";
Trees_din <= "00000110000000000010111101000000";
wait for Clk_period;
Addr <= "0010001000110";
Trees_din <= "00000010000000000100010000100000";
wait for Clk_period;
Addr <= "0010001000111";
Trees_din <= "00000111000000000000101000010000";
wait for Clk_period;
Addr <= "0010001001000";
Trees_din <= "00000001000000000101110000001000";
wait for Clk_period;
Addr <= "0010001001001";
Trees_din <= "00000000000000000011101100000100";
wait for Clk_period;
Addr <= "0010001001010";
Trees_din <= "00000000001000110001001000010001";
wait for Clk_period;
Addr <= "0010001001011";
Trees_din <= "00000000000011110001001000010001";
wait for Clk_period;
Addr <= "0010001001100";
Trees_din <= "00000011000000000011101100000100";
wait for Clk_period;
Addr <= "0010001001101";
Trees_din <= "00000000010001010001001000010001";
wait for Clk_period;
Addr <= "0010001001110";
Trees_din <= "00000000000010110001001000010001";
wait for Clk_period;
Addr <= "0010001001111";
Trees_din <= "00000110000000000010111000001000";
wait for Clk_period;
Addr <= "0010001010000";
Trees_din <= "00000001000000000100100100000100";
wait for Clk_period;
Addr <= "0010001010001";
Trees_din <= "00000000001010000001001000010001";
wait for Clk_period;
Addr <= "0010001010010";
Trees_din <= "00000000010110000001001000010001";
wait for Clk_period;
Addr <= "0010001010011";
Trees_din <= "00000001000000000110000100000100";
wait for Clk_period;
Addr <= "0010001010100";
Trees_din <= "00000000000010110001001000010001";
wait for Clk_period;
Addr <= "0010001010101";
Trees_din <= "00000000010100000001001000010001";
wait for Clk_period;
Addr <= "0010001010110";
Trees_din <= "00000101000000000011101100010000";
wait for Clk_period;
Addr <= "0010001010111";
Trees_din <= "00000000000000000100100100001000";
wait for Clk_period;
Addr <= "0010001011000";
Trees_din <= "00000010000000000101111000000100";
wait for Clk_period;
Addr <= "0010001011001";
Trees_din <= "00000000001011100001001000010001";
wait for Clk_period;
Addr <= "0010001011010";
Trees_din <= "00000000000011010001001000010001";
wait for Clk_period;
Addr <= "0010001011011";
Trees_din <= "00000101000000000000100000000100";
wait for Clk_period;
Addr <= "0010001011100";
Trees_din <= "00000000010110100001001000010001";
wait for Clk_period;
Addr <= "0010001011101";
Trees_din <= "00000000010011000001001000010001";
wait for Clk_period;
Addr <= "0010001011110";
Trees_din <= "00000000000000000110000000001000";
wait for Clk_period;
Addr <= "0010001011111";
Trees_din <= "00000100000000000100101000000100";
wait for Clk_period;
Addr <= "0010001100000";
Trees_din <= "00000000001110100001001000010001";
wait for Clk_period;
Addr <= "0010001100001";
Trees_din <= "00000000001101000001001000010001";
wait for Clk_period;
Addr <= "0010001100010";
Trees_din <= "00000110000000000001010000000100";
wait for Clk_period;
Addr <= "0010001100011";
Trees_din <= "00000000010101110001001000010001";
wait for Clk_period;
Addr <= "0010001100100";
Trees_din <= "00000000000110110001001000010001";
wait for Clk_period;
Addr <= "0010001100101";
Trees_din <= "00000111000000000000001000100000";
wait for Clk_period;
Addr <= "0010001100110";
Trees_din <= "00000111000000000000000000010000";
wait for Clk_period;
Addr <= "0010001100111";
Trees_din <= "00000100000000000010001100001000";
wait for Clk_period;
Addr <= "0010001101000";
Trees_din <= "00000001000000000000110100000100";
wait for Clk_period;
Addr <= "0010001101001";
Trees_din <= "00000000010000000001001000010001";
wait for Clk_period;
Addr <= "0010001101010";
Trees_din <= "00000000010110110001001000010001";
wait for Clk_period;
Addr <= "0010001101011";
Trees_din <= "00000100000000000000000000000100";
wait for Clk_period;
Addr <= "0010001101100";
Trees_din <= "00000000000111110001001000010001";
wait for Clk_period;
Addr <= "0010001101101";
Trees_din <= "00000000010010000001001000010001";
wait for Clk_period;
Addr <= "0010001101110";
Trees_din <= "00000010000000000101111100001000";
wait for Clk_period;
Addr <= "0010001101111";
Trees_din <= "00000110000000000001001100000100";
wait for Clk_period;
Addr <= "0010001110000";
Trees_din <= "00000000010010100001001000010001";
wait for Clk_period;
Addr <= "0010001110001";
Trees_din <= "00000000010111000001001000010001";
wait for Clk_period;
Addr <= "0010001110010";
Trees_din <= "00000010000000000011100000000100";
wait for Clk_period;
Addr <= "0010001110011";
Trees_din <= "00000000011000000001001000010001";
wait for Clk_period;
Addr <= "0010001110100";
Trees_din <= "00000000010111000001001000010001";
wait for Clk_period;
Addr <= "0010001110101";
Trees_din <= "00000001000000000100111100010000";
wait for Clk_period;
Addr <= "0010001110110";
Trees_din <= "00000110000000000100101100001000";
wait for Clk_period;
Addr <= "0010001110111";
Trees_din <= "00000011000000000010110100000100";
wait for Clk_period;
Addr <= "0010001111000";
Trees_din <= "00000000001111110001001000010001";
wait for Clk_period;
Addr <= "0010001111001";
Trees_din <= "00000000011000100001001000010001";
wait for Clk_period;
Addr <= "0010001111010";
Trees_din <= "00000011000000000100110000000100";
wait for Clk_period;
Addr <= "0010001111011";
Trees_din <= "00000000011000110001001000010001";
wait for Clk_period;
Addr <= "0010001111100";
Trees_din <= "00000000010101100001001000010001";
wait for Clk_period;
Addr <= "0010001111101";
Trees_din <= "00000000000000000011011100001000";
wait for Clk_period;
Addr <= "0010001111110";
Trees_din <= "00000100000000000100001000000100";
wait for Clk_period;
Addr <= "0010001111111";
Trees_din <= "00000000001011110001001000010001";
wait for Clk_period;
Addr <= "0010010000000";
Trees_din <= "00000000001000010001001000010001";
wait for Clk_period;
Addr <= "0010010000001";
Trees_din <= "00000011000000000101001100000100";
wait for Clk_period;
Addr <= "0010010000010";
Trees_din <= "00000000001100110001001000010001";
wait for Clk_period;
Addr <= "0010010000011";
Trees_din <= "00000000001011110001001000010001";
wait for Clk_period;



----------tree 9-------------------

Addr <= "0010010000100";
Trees_din <= "00000000000000000100110110000000";
wait for Clk_period;
Addr <= "0010010000101";
Trees_din <= "00000100000000000001110001000000";
wait for Clk_period;
Addr <= "0010010000110";
Trees_din <= "00000011000000000010111000100000";
wait for Clk_period;
Addr <= "0010010000111";
Trees_din <= "00000101000000000011011000010000";
wait for Clk_period;
Addr <= "0010010001000";
Trees_din <= "00000111000000000100011000001000";
wait for Clk_period;
Addr <= "0010010001001";
Trees_din <= "00000000000000000000111000000100";
wait for Clk_period;
Addr <= "0010010001010";
Trees_din <= "00000000011000010001010000001111";
wait for Clk_period;
Addr <= "0010010001011";
Trees_din <= "00000000000001110001010000001111";
wait for Clk_period;
Addr <= "0010010001100";
Trees_din <= "00000010000000000000110000000100";
wait for Clk_period;
Addr <= "0010010001101";
Trees_din <= "00000000000101000001010000001111";
wait for Clk_period;
Addr <= "0010010001110";
Trees_din <= "00000000001101110001010000001111";
wait for Clk_period;
Addr <= "0010010001111";
Trees_din <= "00000001000000000001011000001000";
wait for Clk_period;
Addr <= "0010010010000";
Trees_din <= "00000010000000000101100000000100";
wait for Clk_period;
Addr <= "0010010010001";
Trees_din <= "00000000001001100001010000001111";
wait for Clk_period;
Addr <= "0010010010010";
Trees_din <= "00000000001001000001010000001111";
wait for Clk_period;
Addr <= "0010010010011";
Trees_din <= "00000100000000000010010000000100";
wait for Clk_period;
Addr <= "0010010010100";
Trees_din <= "00000000010011100001010000001111";
wait for Clk_period;
Addr <= "0010010010101";
Trees_din <= "00000000010101110001010000001111";
wait for Clk_period;
Addr <= "0010010010110";
Trees_din <= "00000011000000000000111100010000";
wait for Clk_period;
Addr <= "0010010010111";
Trees_din <= "00000100000000000011100100001000";
wait for Clk_period;
Addr <= "0010010011000";
Trees_din <= "00000011000000000001001000000100";
wait for Clk_period;
Addr <= "0010010011001";
Trees_din <= "00000000001101000001010000001111";
wait for Clk_period;
Addr <= "0010010011010";
Trees_din <= "00000000000010110001010000001111";
wait for Clk_period;
Addr <= "0010010011011";
Trees_din <= "00000101000000000011000000000100";
wait for Clk_period;
Addr <= "0010010011100";
Trees_din <= "00000000001100100001010000001111";
wait for Clk_period;
Addr <= "0010010011101";
Trees_din <= "00000000010100110001010000001111";
wait for Clk_period;
Addr <= "0010010011110";
Trees_din <= "00000011000000000000000000001000";
wait for Clk_period;
Addr <= "0010010011111";
Trees_din <= "00000001000000000001110000000100";
wait for Clk_period;
Addr <= "0010010100000";
Trees_din <= "00000000001101000001010000001111";
wait for Clk_period;
Addr <= "0010010100001";
Trees_din <= "00000000000010010001010000001111";
wait for Clk_period;
Addr <= "0010010100010";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "0010010100011";
Trees_din <= "00000000000101000001010000001111";
wait for Clk_period;
Addr <= "0010010100100";
Trees_din <= "00000000001111100001010000001111";
wait for Clk_period;
Addr <= "0010010100101";
Trees_din <= "00000110000000000001101000100000";
wait for Clk_period;
Addr <= "0010010100110";
Trees_din <= "00000001000000000011111100010000";
wait for Clk_period;
Addr <= "0010010100111";
Trees_din <= "00000101000000000001110000001000";
wait for Clk_period;
Addr <= "0010010101000";
Trees_din <= "00000110000000000001100100000100";
wait for Clk_period;
Addr <= "0010010101001";
Trees_din <= "00000000010000110001010000001111";
wait for Clk_period;
Addr <= "0010010101010";
Trees_din <= "00000000010111000001010000001111";
wait for Clk_period;
Addr <= "0010010101011";
Trees_din <= "00000010000000000001101000000100";
wait for Clk_period;
Addr <= "0010010101100";
Trees_din <= "00000000000001000001010000001111";
wait for Clk_period;
Addr <= "0010010101101";
Trees_din <= "00000000000010000001010000001111";
wait for Clk_period;
Addr <= "0010010101110";
Trees_din <= "00000000000000000011001100001000";
wait for Clk_period;
Addr <= "0010010101111";
Trees_din <= "00000111000000000000011100000100";
wait for Clk_period;
Addr <= "0010010110000";
Trees_din <= "00000000010001110001010000001111";
wait for Clk_period;
Addr <= "0010010110001";
Trees_din <= "00000000010100100001010000001111";
wait for Clk_period;
Addr <= "0010010110010";
Trees_din <= "00000001000000000001100000000100";
wait for Clk_period;
Addr <= "0010010110011";
Trees_din <= "00000000000001110001010000001111";
wait for Clk_period;
Addr <= "0010010110100";
Trees_din <= "00000000000001110001010000001111";
wait for Clk_period;
Addr <= "0010010110101";
Trees_din <= "00000010000000000101111100010000";
wait for Clk_period;
Addr <= "0010010110110";
Trees_din <= "00000110000000000110000100001000";
wait for Clk_period;
Addr <= "0010010110111";
Trees_din <= "00000100000000000010001100000100";
wait for Clk_period;
Addr <= "0010010111000";
Trees_din <= "00000000000011000001010000001111";
wait for Clk_period;
Addr <= "0010010111001";
Trees_din <= "00000000000011100001010000001111";
wait for Clk_period;
Addr <= "0010010111010";
Trees_din <= "00000011000000000101011000000100";
wait for Clk_period;
Addr <= "0010010111011";
Trees_din <= "00000000001111000001010000001111";
wait for Clk_period;
Addr <= "0010010111100";
Trees_din <= "00000000001010110001010000001111";
wait for Clk_period;
Addr <= "0010010111101";
Trees_din <= "00000110000000000001010000001000";
wait for Clk_period;
Addr <= "0010010111110";
Trees_din <= "00000011000000000010110000000100";
wait for Clk_period;
Addr <= "0010010111111";
Trees_din <= "00000000010001110001010000001111";
wait for Clk_period;
Addr <= "0010011000000";
Trees_din <= "00000000000110000001010000001111";
wait for Clk_period;
Addr <= "0010011000001";
Trees_din <= "00000111000000000001001100000100";
wait for Clk_period;
Addr <= "0010011000010";
Trees_din <= "00000000010011010001010000001111";
wait for Clk_period;
Addr <= "0010011000011";
Trees_din <= "00000000010111110001010000001111";
wait for Clk_period;
Addr <= "0010011000100";
Trees_din <= "00000101000000000000111001000000";
wait for Clk_period;
Addr <= "0010011000101";
Trees_din <= "00000011000000000010011000100000";
wait for Clk_period;
Addr <= "0010011000110";
Trees_din <= "00000110000000000100101000010000";
wait for Clk_period;
Addr <= "0010011000111";
Trees_din <= "00000100000000000011110100001000";
wait for Clk_period;
Addr <= "0010011001000";
Trees_din <= "00000011000000000100010100000100";
wait for Clk_period;
Addr <= "0010011001001";
Trees_din <= "00000000001110100001010000001111";
wait for Clk_period;
Addr <= "0010011001010";
Trees_din <= "00000000000010100001010000001111";
wait for Clk_period;
Addr <= "0010011001011";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "0010011001100";
Trees_din <= "00000000001001010001010000001111";
wait for Clk_period;
Addr <= "0010011001101";
Trees_din <= "00000000001001100001010000001111";
wait for Clk_period;
Addr <= "0010011001110";
Trees_din <= "00000101000000000101001100001000";
wait for Clk_period;
Addr <= "0010011001111";
Trees_din <= "00000011000000000010111100000100";
wait for Clk_period;
Addr <= "0010011010000";
Trees_din <= "00000000001000100001010000001111";
wait for Clk_period;
Addr <= "0010011010001";
Trees_din <= "00000000010010000001010000001111";
wait for Clk_period;
Addr <= "0010011010010";
Trees_din <= "00000111000000000000100100000100";
wait for Clk_period;
Addr <= "0010011010011";
Trees_din <= "00000000000000010001010000001111";
wait for Clk_period;
Addr <= "0010011010100";
Trees_din <= "00000000000111010001010000001111";
wait for Clk_period;
Addr <= "0010011010101";
Trees_din <= "00000001000000000000000100010000";
wait for Clk_period;
Addr <= "0010011010110";
Trees_din <= "00000011000000000101010000001000";
wait for Clk_period;
Addr <= "0010011010111";
Trees_din <= "00000110000000000100010100000100";
wait for Clk_period;
Addr <= "0010011011000";
Trees_din <= "00000000010101010001010000001111";
wait for Clk_period;
Addr <= "0010011011001";
Trees_din <= "00000000010110000001010000001111";
wait for Clk_period;
Addr <= "0010011011010";
Trees_din <= "00000010000000000101010100000100";
wait for Clk_period;
Addr <= "0010011011011";
Trees_din <= "00000000001110100001010000001111";
wait for Clk_period;
Addr <= "0010011011100";
Trees_din <= "00000000000101000001010000001111";
wait for Clk_period;
Addr <= "0010011011101";
Trees_din <= "00000100000000000110000100001000";
wait for Clk_period;
Addr <= "0010011011110";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "0010011011111";
Trees_din <= "00000000001111110001010000001111";
wait for Clk_period;
Addr <= "0010011100000";
Trees_din <= "00000000010011010001010000001111";
wait for Clk_period;
Addr <= "0010011100001";
Trees_din <= "00000101000000000011000100000100";
wait for Clk_period;
Addr <= "0010011100010";
Trees_din <= "00000000010100100001010000001111";
wait for Clk_period;
Addr <= "0010011100011";
Trees_din <= "00000000000000000001010000001111";
wait for Clk_period;
Addr <= "0010011100100";
Trees_din <= "00000100000000000011001100100000";
wait for Clk_period;
Addr <= "0010011100101";
Trees_din <= "00000000000000000101010000010000";
wait for Clk_period;
Addr <= "0010011100110";
Trees_din <= "00000011000000000011011000001000";
wait for Clk_period;
Addr <= "0010011100111";
Trees_din <= "00000100000000000010111000000100";
wait for Clk_period;
Addr <= "0010011101000";
Trees_din <= "00000000010110010001010000001111";
wait for Clk_period;
Addr <= "0010011101001";
Trees_din <= "00000000000001010001010000001111";
wait for Clk_period;
Addr <= "0010011101010";
Trees_din <= "00000111000000000000111000000100";
wait for Clk_period;
Addr <= "0010011101011";
Trees_din <= "00000000010011100001010000001111";
wait for Clk_period;
Addr <= "0010011101100";
Trees_din <= "00000000010000010001010000001111";
wait for Clk_period;
Addr <= "0010011101101";
Trees_din <= "00000111000000000001111000001000";
wait for Clk_period;
Addr <= "0010011101110";
Trees_din <= "00000000000000000011001100000100";
wait for Clk_period;
Addr <= "0010011101111";
Trees_din <= "00000000010111100001010000001111";
wait for Clk_period;
Addr <= "0010011110000";
Trees_din <= "00000000010101110001010000001111";
wait for Clk_period;
Addr <= "0010011110001";
Trees_din <= "00000011000000000100011100000100";
wait for Clk_period;
Addr <= "0010011110010";
Trees_din <= "00000000010001000001010000001111";
wait for Clk_period;
Addr <= "0010011110011";
Trees_din <= "00000000010111010001010000001111";
wait for Clk_period;
Addr <= "0010011110100";
Trees_din <= "00000111000000000101001000010000";
wait for Clk_period;
Addr <= "0010011110101";
Trees_din <= "00000110000000000000110000001000";
wait for Clk_period;
Addr <= "0010011110110";
Trees_din <= "00000011000000000000101000000100";
wait for Clk_period;
Addr <= "0010011110111";
Trees_din <= "00000000010111010001010000001111";
wait for Clk_period;
Addr <= "0010011111000";
Trees_din <= "00000000010001110001010000001111";
wait for Clk_period;
Addr <= "0010011111001";
Trees_din <= "00000011000000000100000000000100";
wait for Clk_period;
Addr <= "0010011111010";
Trees_din <= "00000000000000110001010000001111";
wait for Clk_period;
Addr <= "0010011111011";
Trees_din <= "00000000001000000001010000001111";
wait for Clk_period;
Addr <= "0010011111100";
Trees_din <= "00000000000000000101100000001000";
wait for Clk_period;
Addr <= "0010011111101";
Trees_din <= "00000110000000000110001100000100";
wait for Clk_period;
Addr <= "0010011111110";
Trees_din <= "00000000001110010001010000001111";
wait for Clk_period;
Addr <= "0010011111111";
Trees_din <= "00000000000101000001010000001111";
wait for Clk_period;
Addr <= "0010100000000";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "0010100000001";
Trees_din <= "00000000001100110001010000001111";
wait for Clk_period;
Addr <= "0010100000010";
Trees_din <= "00000000000101100001010000001111";
wait for Clk_period;



----------tree 10-------------------

Addr <= "0010100000011";
Trees_din <= "00000100000000000001111110000000";
wait for Clk_period;
Addr <= "0010100000100";
Trees_din <= "00000111000000000000010101000000";
wait for Clk_period;
Addr <= "0010100000101";
Trees_din <= "00000000000000000100000100100000";
wait for Clk_period;
Addr <= "0010100000110";
Trees_din <= "00000000000000000011011100010000";
wait for Clk_period;
Addr <= "0010100000111";
Trees_din <= "00000001000000000001011000001000";
wait for Clk_period;
Addr <= "0010100001000";
Trees_din <= "00000011000000000011110100000100";
wait for Clk_period;
Addr <= "0010100001001";
Trees_din <= "00000000001110110001011000001001";
wait for Clk_period;
Addr <= "0010100001010";
Trees_din <= "00000000000011000001011000001001";
wait for Clk_period;
Addr <= "0010100001011";
Trees_din <= "00000111000000000010011000000100";
wait for Clk_period;
Addr <= "0010100001100";
Trees_din <= "00000000000111010001011000001001";
wait for Clk_period;
Addr <= "0010100001101";
Trees_din <= "00000000010000010001011000001001";
wait for Clk_period;
Addr <= "0010100001110";
Trees_din <= "00000011000000000011100000001000";
wait for Clk_period;
Addr <= "0010100001111";
Trees_din <= "00000101000000000101101100000100";
wait for Clk_period;
Addr <= "0010100010000";
Trees_din <= "00000000001101110001011000001001";
wait for Clk_period;
Addr <= "0010100010001";
Trees_din <= "00000000000100000001011000001001";
wait for Clk_period;
Addr <= "0010100010010";
Trees_din <= "00000000000000000011001100000100";
wait for Clk_period;
Addr <= "0010100010011";
Trees_din <= "00000000001001110001011000001001";
wait for Clk_period;
Addr <= "0010100010100";
Trees_din <= "00000000000100110001011000001001";
wait for Clk_period;
Addr <= "0010100010101";
Trees_din <= "00000100000000000001111000010000";
wait for Clk_period;
Addr <= "0010100010110";
Trees_din <= "00000101000000000011100100001000";
wait for Clk_period;
Addr <= "0010100010111";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "0010100011000";
Trees_din <= "00000000001000000001011000001001";
wait for Clk_period;
Addr <= "0010100011001";
Trees_din <= "00000000000001000001011000001001";
wait for Clk_period;
Addr <= "0010100011010";
Trees_din <= "00000100000000000001100000000100";
wait for Clk_period;
Addr <= "0010100011011";
Trees_din <= "00000000000010000001011000001001";
wait for Clk_period;
Addr <= "0010100011100";
Trees_din <= "00000000010111110001011000001001";
wait for Clk_period;
Addr <= "0010100011101";
Trees_din <= "00000000000000000101111000001000";
wait for Clk_period;
Addr <= "0010100011110";
Trees_din <= "00000011000000000000011100000100";
wait for Clk_period;
Addr <= "0010100011111";
Trees_din <= "00000000010100000001011000001001";
wait for Clk_period;
Addr <= "0010100100000";
Trees_din <= "00000000001001110001011000001001";
wait for Clk_period;
Addr <= "0010100100001";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0010100100010";
Trees_din <= "00000000010010000001011000001001";
wait for Clk_period;
Addr <= "0010100100011";
Trees_din <= "00000000001111100001011000001001";
wait for Clk_period;
Addr <= "0010100100100";
Trees_din <= "00000101000000000101000000100000";
wait for Clk_period;
Addr <= "0010100100101";
Trees_din <= "00000100000000000000101100010000";
wait for Clk_period;
Addr <= "0010100100110";
Trees_din <= "00000001000000000000101000001000";
wait for Clk_period;
Addr <= "0010100100111";
Trees_din <= "00000100000000000001011100000100";
wait for Clk_period;
Addr <= "0010100101000";
Trees_din <= "00000000010110000001011000001001";
wait for Clk_period;
Addr <= "0010100101001";
Trees_din <= "00000000000111100001011000001001";
wait for Clk_period;
Addr <= "0010100101010";
Trees_din <= "00000111000000000000110100000100";
wait for Clk_period;
Addr <= "0010100101011";
Trees_din <= "00000000000011000001011000001001";
wait for Clk_period;
Addr <= "0010100101100";
Trees_din <= "00000000000101000001011000001001";
wait for Clk_period;
Addr <= "0010100101101";
Trees_din <= "00000111000000000110010000001000";
wait for Clk_period;
Addr <= "0010100101110";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "0010100101111";
Trees_din <= "00000000010110110001011000001001";
wait for Clk_period;
Addr <= "0010100110000";
Trees_din <= "00000000001111000001011000001001";
wait for Clk_period;
Addr <= "0010100110001";
Trees_din <= "00000000000000000101101100000100";
wait for Clk_period;
Addr <= "0010100110010";
Trees_din <= "00000000010001010001011000001001";
wait for Clk_period;
Addr <= "0010100110011";
Trees_din <= "00000000010101110001011000001001";
wait for Clk_period;
Addr <= "0010100110100";
Trees_din <= "00000001000000000000100000010000";
wait for Clk_period;
Addr <= "0010100110101";
Trees_din <= "00000001000000000000011100001000";
wait for Clk_period;
Addr <= "0010100110110";
Trees_din <= "00000101000000000110001100000100";
wait for Clk_period;
Addr <= "0010100110111";
Trees_din <= "00000000010101000001011000001001";
wait for Clk_period;
Addr <= "0010100111000";
Trees_din <= "00000000001010110001011000001001";
wait for Clk_period;
Addr <= "0010100111001";
Trees_din <= "00000010000000000100010000000100";
wait for Clk_period;
Addr <= "0010100111010";
Trees_din <= "00000000001001100001011000001001";
wait for Clk_period;
Addr <= "0010100111011";
Trees_din <= "00000000000001010001011000001001";
wait for Clk_period;
Addr <= "0010100111100";
Trees_din <= "00000110000000000011010100001000";
wait for Clk_period;
Addr <= "0010100111101";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0010100111110";
Trees_din <= "00000000001101010001011000001001";
wait for Clk_period;
Addr <= "0010100111111";
Trees_din <= "00000000000001010001011000001001";
wait for Clk_period;
Addr <= "0010101000000";
Trees_din <= "00000101000000000000000000000100";
wait for Clk_period;
Addr <= "0010101000001";
Trees_din <= "00000000010100000001011000001001";
wait for Clk_period;
Addr <= "0010101000010";
Trees_din <= "00000000001001110001011000001001";
wait for Clk_period;
Addr <= "0010101000011";
Trees_din <= "00000011000000000011100101000000";
wait for Clk_period;
Addr <= "0010101000100";
Trees_din <= "00000110000000000011011000100000";
wait for Clk_period;
Addr <= "0010101000101";
Trees_din <= "00000010000000000101001100010000";
wait for Clk_period;
Addr <= "0010101000110";
Trees_din <= "00000110000000000010100000001000";
wait for Clk_period;
Addr <= "0010101000111";
Trees_din <= "00000110000000000001001000000100";
wait for Clk_period;
Addr <= "0010101001000";
Trees_din <= "00000000000100000001011000001001";
wait for Clk_period;
Addr <= "0010101001001";
Trees_din <= "00000000001100110001011000001001";
wait for Clk_period;
Addr <= "0010101001010";
Trees_din <= "00000010000000000000000000000100";
wait for Clk_period;
Addr <= "0010101001011";
Trees_din <= "00000000001011100001011000001001";
wait for Clk_period;
Addr <= "0010101001100";
Trees_din <= "00000000001011010001011000001001";
wait for Clk_period;
Addr <= "0010101001101";
Trees_din <= "00000011000000000010111000001000";
wait for Clk_period;
Addr <= "0010101001110";
Trees_din <= "00000001000000000001110000000100";
wait for Clk_period;
Addr <= "0010101001111";
Trees_din <= "00000000001110100001011000001001";
wait for Clk_period;
Addr <= "0010101010000";
Trees_din <= "00000000011000100001011000001001";
wait for Clk_period;
Addr <= "0010101010001";
Trees_din <= "00000101000000000100110100000100";
wait for Clk_period;
Addr <= "0010101010010";
Trees_din <= "00000000001111000001011000001001";
wait for Clk_period;
Addr <= "0010101010011";
Trees_din <= "00000000000000110001011000001001";
wait for Clk_period;
Addr <= "0010101010100";
Trees_din <= "00000101000000000000001100010000";
wait for Clk_period;
Addr <= "0010101010101";
Trees_din <= "00000111000000000010110100001000";
wait for Clk_period;
Addr <= "0010101010110";
Trees_din <= "00000100000000000101100100000100";
wait for Clk_period;
Addr <= "0010101010111";
Trees_din <= "00000000001010000001011000001001";
wait for Clk_period;
Addr <= "0010101011000";
Trees_din <= "00000000001101010001011000001001";
wait for Clk_period;
Addr <= "0010101011001";
Trees_din <= "00000101000000000110001000000100";
wait for Clk_period;
Addr <= "0010101011010";
Trees_din <= "00000000010101110001011000001001";
wait for Clk_period;
Addr <= "0010101011011";
Trees_din <= "00000000000101100001011000001001";
wait for Clk_period;
Addr <= "0010101011100";
Trees_din <= "00000010000000000100110000001000";
wait for Clk_period;
Addr <= "0010101011101";
Trees_din <= "00000110000000000011110000000100";
wait for Clk_period;
Addr <= "0010101011110";
Trees_din <= "00000000010101010001011000001001";
wait for Clk_period;
Addr <= "0010101011111";
Trees_din <= "00000000001001110001011000001001";
wait for Clk_period;
Addr <= "0010101100000";
Trees_din <= "00000101000000000011001000000100";
wait for Clk_period;
Addr <= "0010101100001";
Trees_din <= "00000000000000110001011000001001";
wait for Clk_period;
Addr <= "0010101100010";
Trees_din <= "00000000001101110001011000001001";
wait for Clk_period;
Addr <= "0010101100011";
Trees_din <= "00000010000000000011110100100000";
wait for Clk_period;
Addr <= "0010101100100";
Trees_din <= "00000001000000000010011000010000";
wait for Clk_period;
Addr <= "0010101100101";
Trees_din <= "00000010000000000001101100001000";
wait for Clk_period;
Addr <= "0010101100110";
Trees_din <= "00000011000000000011101000000100";
wait for Clk_period;
Addr <= "0010101100111";
Trees_din <= "00000000001110010001011000001001";
wait for Clk_period;
Addr <= "0010101101000";
Trees_din <= "00000000001010000001011000001001";
wait for Clk_period;
Addr <= "0010101101001";
Trees_din <= "00000111000000000100000100000100";
wait for Clk_period;
Addr <= "0010101101010";
Trees_din <= "00000000001100010001011000001001";
wait for Clk_period;
Addr <= "0010101101011";
Trees_din <= "00000000010111110001011000001001";
wait for Clk_period;
Addr <= "0010101101100";
Trees_din <= "00000011000000000000110000001000";
wait for Clk_period;
Addr <= "0010101101101";
Trees_din <= "00000101000000000000111000000100";
wait for Clk_period;
Addr <= "0010101101110";
Trees_din <= "00000000010101110001011000001001";
wait for Clk_period;
Addr <= "0010101101111";
Trees_din <= "00000000001000000001011000001001";
wait for Clk_period;
Addr <= "0010101110000";
Trees_din <= "00000110000000000010000100000100";
wait for Clk_period;
Addr <= "0010101110001";
Trees_din <= "00000000001011000001011000001001";
wait for Clk_period;
Addr <= "0010101110010";
Trees_din <= "00000000000110010001011000001001";
wait for Clk_period;
Addr <= "0010101110011";
Trees_din <= "00000111000000000101101000010000";
wait for Clk_period;
Addr <= "0010101110100";
Trees_din <= "00000111000000000011011100001000";
wait for Clk_period;
Addr <= "0010101110101";
Trees_din <= "00000010000000000101011100000100";
wait for Clk_period;
Addr <= "0010101110110";
Trees_din <= "00000000000101100001011000001001";
wait for Clk_period;
Addr <= "0010101110111";
Trees_din <= "00000000000101010001011000001001";
wait for Clk_period;
Addr <= "0010101111000";
Trees_din <= "00000111000000000000100000000100";
wait for Clk_period;
Addr <= "0010101111001";
Trees_din <= "00000000000000110001011000001001";
wait for Clk_period;
Addr <= "0010101111010";
Trees_din <= "00000000000111010001011000001001";
wait for Clk_period;
Addr <= "0010101111011";
Trees_din <= "00000010000000000011001000001000";
wait for Clk_period;
Addr <= "0010101111100";
Trees_din <= "00000011000000000011011100000100";
wait for Clk_period;
Addr <= "0010101111101";
Trees_din <= "00000000001011010001011000001001";
wait for Clk_period;
Addr <= "0010101111110";
Trees_din <= "00000000010000000001011000001001";
wait for Clk_period;
Addr <= "0010101111111";
Trees_din <= "00000010000000000010101100000100";
wait for Clk_period;
Addr <= "0010110000000";
Trees_din <= "00000000001011000001011000001001";
wait for Clk_period;
Addr <= "0010110000001";
Trees_din <= "00000000001111010001011000001001";
wait for Clk_period;



----------tree 11-------------------

Addr <= "0010110000010";
Trees_din <= "00000011000000000101000110000000";
wait for Clk_period;
Addr <= "0010110000011";
Trees_din <= "00000110000000000010000101000000";
wait for Clk_period;
Addr <= "0010110000100";
Trees_din <= "00000000000000000010110100100000";
wait for Clk_period;
Addr <= "0010110000101";
Trees_din <= "00000001000000000001110000010000";
wait for Clk_period;
Addr <= "0010110000110";
Trees_din <= "00000111000000000011101100001000";
wait for Clk_period;
Addr <= "0010110000111";
Trees_din <= "00000101000000000001010000000100";
wait for Clk_period;
Addr <= "0010110001000";
Trees_din <= "00000000001010100000000000000011";
wait for Clk_period;
Addr <= "0010110001001";
Trees_din <= "00000000010011110000000000000011";
wait for Clk_period;
Addr <= "0010110001010";
Trees_din <= "00000001000000000000110100000100";
wait for Clk_period;
Addr <= "0010110001011";
Trees_din <= "00000000010011000000000000000011";
wait for Clk_period;
Addr <= "0010110001100";
Trees_din <= "00000000010110110000000000000011";
wait for Clk_period;
Addr <= "0010110001101";
Trees_din <= "00000110000000000110001000001000";
wait for Clk_period;
Addr <= "0010110001110";
Trees_din <= "00000011000000000011011000000100";
wait for Clk_period;
Addr <= "0010110001111";
Trees_din <= "00000000011001000000000000000011";
wait for Clk_period;
Addr <= "0010110010000";
Trees_din <= "00000000000110000000000000000011";
wait for Clk_period;
Addr <= "0010110010001";
Trees_din <= "00000100000000000110010000000100";
wait for Clk_period;
Addr <= "0010110010010";
Trees_din <= "00000000010011110000000000000011";
wait for Clk_period;
Addr <= "0010110010011";
Trees_din <= "00000000000000010000000000000011";
wait for Clk_period;
Addr <= "0010110010100";
Trees_din <= "00000001000000000100010100010000";
wait for Clk_period;
Addr <= "0010110010101";
Trees_din <= "00000011000000000010000000001000";
wait for Clk_period;
Addr <= "0010110010110";
Trees_din <= "00000100000000000101101100000100";
wait for Clk_period;
Addr <= "0010110010111";
Trees_din <= "00000000010011010000000000000011";
wait for Clk_period;
Addr <= "0010110011000";
Trees_din <= "00000000001110000000000000000011";
wait for Clk_period;
Addr <= "0010110011001";
Trees_din <= "00000010000000000011111100000100";
wait for Clk_period;
Addr <= "0010110011010";
Trees_din <= "00000000010010010000000000000011";
wait for Clk_period;
Addr <= "0010110011011";
Trees_din <= "00000000001001110000000000000011";
wait for Clk_period;
Addr <= "0010110011100";
Trees_din <= "00000011000000000100100000001000";
wait for Clk_period;
Addr <= "0010110011101";
Trees_din <= "00000111000000000011111100000100";
wait for Clk_period;
Addr <= "0010110011110";
Trees_din <= "00000000001110000000000000000011";
wait for Clk_period;
Addr <= "0010110011111";
Trees_din <= "00000000010010010000000000000011";
wait for Clk_period;
Addr <= "0010110100000";
Trees_din <= "00000010000000000000101100000100";
wait for Clk_period;
Addr <= "0010110100001";
Trees_din <= "00000000000010100000000000000011";
wait for Clk_period;
Addr <= "0010110100010";
Trees_din <= "00000000010000110000000000000011";
wait for Clk_period;
Addr <= "0010110100011";
Trees_din <= "00000110000000000101010100100000";
wait for Clk_period;
Addr <= "0010110100100";
Trees_din <= "00000001000000000000010000010000";
wait for Clk_period;
Addr <= "0010110100101";
Trees_din <= "00000100000000000100110000001000";
wait for Clk_period;
Addr <= "0010110100110";
Trees_din <= "00000100000000000001110100000100";
wait for Clk_period;
Addr <= "0010110100111";
Trees_din <= "00000000011000110000000000000011";
wait for Clk_period;
Addr <= "0010110101000";
Trees_din <= "00000000010001100000000000000011";
wait for Clk_period;
Addr <= "0010110101001";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0010110101010";
Trees_din <= "00000000001011000000000000000011";
wait for Clk_period;
Addr <= "0010110101011";
Trees_din <= "00000000000110100000000000000011";
wait for Clk_period;
Addr <= "0010110101100";
Trees_din <= "00000010000000000100000000001000";
wait for Clk_period;
Addr <= "0010110101101";
Trees_din <= "00000011000000000010010000000100";
wait for Clk_period;
Addr <= "0010110101110";
Trees_din <= "00000000000011000000000000000011";
wait for Clk_period;
Addr <= "0010110101111";
Trees_din <= "00000000000010100000000000000011";
wait for Clk_period;
Addr <= "0010110110000";
Trees_din <= "00000101000000000000111100000100";
wait for Clk_period;
Addr <= "0010110110001";
Trees_din <= "00000000001011010000000000000011";
wait for Clk_period;
Addr <= "0010110110010";
Trees_din <= "00000000010001010000000000000011";
wait for Clk_period;
Addr <= "0010110110011";
Trees_din <= "00000000000000000011110000010000";
wait for Clk_period;
Addr <= "0010110110100";
Trees_din <= "00000010000000000101111000001000";
wait for Clk_period;
Addr <= "0010110110101";
Trees_din <= "00000111000000000100101100000100";
wait for Clk_period;
Addr <= "0010110110110";
Trees_din <= "00000000000110100000000000000011";
wait for Clk_period;
Addr <= "0010110110111";
Trees_din <= "00000000001011010000000000000011";
wait for Clk_period;
Addr <= "0010110111000";
Trees_din <= "00000011000000000000111000000100";
wait for Clk_period;
Addr <= "0010110111001";
Trees_din <= "00000000000101110000000000000011";
wait for Clk_period;
Addr <= "0010110111010";
Trees_din <= "00000000010101100000000000000011";
wait for Clk_period;
Addr <= "0010110111011";
Trees_din <= "00000111000000000011000100001000";
wait for Clk_period;
Addr <= "0010110111100";
Trees_din <= "00000010000000000000110100000100";
wait for Clk_period;
Addr <= "0010110111101";
Trees_din <= "00000000000100000000000000000011";
wait for Clk_period;
Addr <= "0010110111110";
Trees_din <= "00000000010101000000000000000011";
wait for Clk_period;
Addr <= "0010110111111";
Trees_din <= "00000101000000000100001100000100";
wait for Clk_period;
Addr <= "0010111000000";
Trees_din <= "00000000000000110000000000000011";
wait for Clk_period;
Addr <= "0010111000001";
Trees_din <= "00000000001010100000000000000011";
wait for Clk_period;
Addr <= "0010111000010";
Trees_din <= "00000000000000000100100001000000";
wait for Clk_period;
Addr <= "0010111000011";
Trees_din <= "00000101000000000000101100100000";
wait for Clk_period;
Addr <= "0010111000100";
Trees_din <= "00000010000000000010111100010000";
wait for Clk_period;
Addr <= "0010111000101";
Trees_din <= "00000011000000000010111100001000";
wait for Clk_period;
Addr <= "0010111000110";
Trees_din <= "00000010000000000001110000000100";
wait for Clk_period;
Addr <= "0010111000111";
Trees_din <= "00000000010011110000000000000011";
wait for Clk_period;
Addr <= "0010111001000";
Trees_din <= "00000000000000100000000000000011";
wait for Clk_period;
Addr <= "0010111001001";
Trees_din <= "00000010000000000011011100000100";
wait for Clk_period;
Addr <= "0010111001010";
Trees_din <= "00000000000001100000000000000011";
wait for Clk_period;
Addr <= "0010111001011";
Trees_din <= "00000000000101000000000000000011";
wait for Clk_period;
Addr <= "0010111001100";
Trees_din <= "00000010000000000000101100001000";
wait for Clk_period;
Addr <= "0010111001101";
Trees_din <= "00000000000000000000001100000100";
wait for Clk_period;
Addr <= "0010111001110";
Trees_din <= "00000000010010000000000000000011";
wait for Clk_period;
Addr <= "0010111001111";
Trees_din <= "00000000010111110000000000000011";
wait for Clk_period;
Addr <= "0010111010000";
Trees_din <= "00000100000000000010110100000100";
wait for Clk_period;
Addr <= "0010111010001";
Trees_din <= "00000000000100010000000000000011";
wait for Clk_period;
Addr <= "0010111010010";
Trees_din <= "00000000000011110000000000000011";
wait for Clk_period;
Addr <= "0010111010011";
Trees_din <= "00000001000000000101001000010000";
wait for Clk_period;
Addr <= "0010111010100";
Trees_din <= "00000101000000000101010100001000";
wait for Clk_period;
Addr <= "0010111010101";
Trees_din <= "00000100000000000100001100000100";
wait for Clk_period;
Addr <= "0010111010110";
Trees_din <= "00000000000011010000000000000011";
wait for Clk_period;
Addr <= "0010111010111";
Trees_din <= "00000000000110010000000000000011";
wait for Clk_period;
Addr <= "0010111011000";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "0010111011001";
Trees_din <= "00000000010000000000000000000011";
wait for Clk_period;
Addr <= "0010111011010";
Trees_din <= "00000000010011110000000000000011";
wait for Clk_period;
Addr <= "0010111011011";
Trees_din <= "00000001000000000101000000001000";
wait for Clk_period;
Addr <= "0010111011100";
Trees_din <= "00000101000000000000011000000100";
wait for Clk_period;
Addr <= "0010111011101";
Trees_din <= "00000000001010010000000000000011";
wait for Clk_period;
Addr <= "0010111011110";
Trees_din <= "00000000000000000000000000000011";
wait for Clk_period;
Addr <= "0010111011111";
Trees_din <= "00000001000000000101000100000100";
wait for Clk_period;
Addr <= "0010111100000";
Trees_din <= "00000000000100110000000000000011";
wait for Clk_period;
Addr <= "0010111100001";
Trees_din <= "00000000000001010000000000000011";
wait for Clk_period;
Addr <= "0010111100010";
Trees_din <= "00000010000000000010100000100000";
wait for Clk_period;
Addr <= "0010111100011";
Trees_din <= "00000001000000000011100100010000";
wait for Clk_period;
Addr <= "0010111100100";
Trees_din <= "00000000000000000100000000001000";
wait for Clk_period;
Addr <= "0010111100101";
Trees_din <= "00000111000000000000110100000100";
wait for Clk_period;
Addr <= "0010111100110";
Trees_din <= "00000000001111110000000000000011";
wait for Clk_period;
Addr <= "0010111100111";
Trees_din <= "00000000000001100000000000000011";
wait for Clk_period;
Addr <= "0010111101000";
Trees_din <= "00000100000000000010001100000100";
wait for Clk_period;
Addr <= "0010111101001";
Trees_din <= "00000000010110100000000000000011";
wait for Clk_period;
Addr <= "0010111101010";
Trees_din <= "00000000010110100000000000000011";
wait for Clk_period;
Addr <= "0010111101011";
Trees_din <= "00000110000000000101100100001000";
wait for Clk_period;
Addr <= "0010111101100";
Trees_din <= "00000001000000000011011100000100";
wait for Clk_period;
Addr <= "0010111101101";
Trees_din <= "00000000000011100000000000000011";
wait for Clk_period;
Addr <= "0010111101110";
Trees_din <= "00000000010010100000000000000011";
wait for Clk_period;
Addr <= "0010111101111";
Trees_din <= "00000000000000000000010000000100";
wait for Clk_period;
Addr <= "0010111110000";
Trees_din <= "00000000010010100000000000000011";
wait for Clk_period;
Addr <= "0010111110001";
Trees_din <= "00000000000001010000000000000011";
wait for Clk_period;
Addr <= "0010111110010";
Trees_din <= "00000111000000000100100100010000";
wait for Clk_period;
Addr <= "0010111110011";
Trees_din <= "00000011000000000011000000001000";
wait for Clk_period;
Addr <= "0010111110100";
Trees_din <= "00000111000000000000010000000100";
wait for Clk_period;
Addr <= "0010111110101";
Trees_din <= "00000000001001110000000000000011";
wait for Clk_period;
Addr <= "0010111110110";
Trees_din <= "00000000010100100000000000000011";
wait for Clk_period;
Addr <= "0010111110111";
Trees_din <= "00000111000000000000011100000100";
wait for Clk_period;
Addr <= "0010111111000";
Trees_din <= "00000000000111110000000000000011";
wait for Clk_period;
Addr <= "0010111111001";
Trees_din <= "00000000000110010000000000000011";
wait for Clk_period;
Addr <= "0010111111010";
Trees_din <= "00000110000000000000010000001000";
wait for Clk_period;
Addr <= "0010111111011";
Trees_din <= "00000111000000000011000100000100";
wait for Clk_period;
Addr <= "0010111111100";
Trees_din <= "00000000011001000000000000000011";
wait for Clk_period;
Addr <= "0010111111101";
Trees_din <= "00000000010110110000000000000011";
wait for Clk_period;
Addr <= "0010111111110";
Trees_din <= "00000001000000000011011100000100";
wait for Clk_period;
Addr <= "0010111111111";
Trees_din <= "00000000000001110000000000000011";
wait for Clk_period;
Addr <= "0011000000000";
Trees_din <= "00000000000000100000000000000011";
wait for Clk_period;


-- LOAD TREES END
-----------------------------------------------------------------------

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period;

        -- class_label <= std_logic_vector(to_unsigned(0, class_label'length));

        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';

-- LOAD FEATURES START
-----------------------------------------------------------------------

        Features_din <= "0000000000110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';

        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;

        Last_feature <= '1';
        pc_count     <= '1';
        Features_din <= "0000000000110010";
        wait for Clk_period;

-- LOAD FEATURES START
-----------------------------------------------------------------------

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';

        -- Wait until inference is complete
        v_TIME := now;
        wait until Finish = '1';
        v_TIME := now - V_TIME;
        report "Execution Time = " & time'image(v_TIME);

        wait for Clk_period * 1/2;

        if Dout = class_label then
            hc_count <= '1';
        end if;

        wait for Clk_period;
        hc_count <= '0';

        stop;
    end process;
end;
    