
-------------------------------------------------------------------------------
-- VHDL test file for 'image.vhd'
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;
use std.env.stop;

entity image_test is
    generic(TREE_RAM_BITS: positive := 13;
            NUM_CLASSES:   positive := 2;
            NUM_FEATURES:  positive := 8);
end image_test;

architecture behavior of image_test is

    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;

             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);

             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;

             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;

    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;

    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto 0);
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';

    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);

    -- Clock period definition
    constant Clk_period : time := 10 ns;

    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');

    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

    -------------------- Newly added signals --------------------

    -- signal addr_count, addr_count_n: std_logic_vector(TREE_RAM_BITS - 1 downto 0);
    shared variable v_TIME : time := 0 ns;

begin

    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);

    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);

    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);

    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;

    -- Stimulus process
    stim_proc: process
    begin

        Reset <= '1';
        Addr <= "0000000000000";

        -- hold reset state for 100 ns.
        wait for 100 ns;

        Reset <= '0';

        wait for Clk_period*10;


-- LOAD TREES START
-----------------------------------------------------------------------

-- Class number = 2
-- Max depth = 7
-- Min depth = 7
-- Tree number = 60
-- average stand deviation for each class is: 
-- class 0 = 0.0
-- class 1 = 0.0

-- LOAD TREES
-----------------------------------------------------------------------

-- Load and valid trees flags
Load_trees <= '1';
Valid_node <= '1';

-- load tree numbers 
Addr <= "0000000000000";
Trees_din <= x"0000003c";
wait for Clk_period;

-- Reset load flag
Load_trees <= '0';    
    
-- Load starting address
--tree 0 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000001";
Trees_din <= "00000000000000000000000000111101";
wait for Clk_period;

--tree 1 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000010";
Trees_din <= "00000000000000000000000010111100";
wait for Clk_period;

--tree 2 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000011";
Trees_din <= "00000000000000000000000100111011";
wait for Clk_period;

--tree 3 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000100";
Trees_din <= "00000000000000000000000110111010";
wait for Clk_period;

--tree 4 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000101";
Trees_din <= "00000000000000000000001000111001";
wait for Clk_period;

--tree 5 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000110";
Trees_din <= "00000000000000000000001010111000";
wait for Clk_period;

--tree 6 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000000111";
Trees_din <= "00000000000000000000001100110111";
wait for Clk_period;

--tree 7 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001000";
Trees_din <= "00000000000000000000001110110110";
wait for Clk_period;

--tree 8 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001001";
Trees_din <= "00000000000000000000010000110101";
wait for Clk_period;

--tree 9 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001010";
Trees_din <= "00000000000000000000010010110100";
wait for Clk_period;

--tree 10 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001011";
Trees_din <= "00000000000000000000010100110011";
wait for Clk_period;

--tree 11 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001100";
Trees_din <= "00000000000000000000010110110010";
wait for Clk_period;

--tree 12 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001101";
Trees_din <= "00000000000000000000011000110001";
wait for Clk_period;

--tree 13 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001110";
Trees_din <= "00000000000000000000011010110000";
wait for Clk_period;

--tree 14 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000001111";
Trees_din <= "00000000000000000000011100101111";
wait for Clk_period;

--tree 15 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010000";
Trees_din <= "00000000000000000000011110101110";
wait for Clk_period;

--tree 16 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010001";
Trees_din <= "00000000000000000000100000101101";
wait for Clk_period;

--tree 17 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010010";
Trees_din <= "00000000000000000000100010101100";
wait for Clk_period;

--tree 18 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010011";
Trees_din <= "00000000000000000000100100101011";
wait for Clk_period;

--tree 19 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010100";
Trees_din <= "00000000000000000000100110101010";
wait for Clk_period;

--tree 20 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010101";
Trees_din <= "00000000000000000000101000101001";
wait for Clk_period;

--tree 21 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010110";
Trees_din <= "00000000000000000000101010101000";
wait for Clk_period;

--tree 22 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000010111";
Trees_din <= "00000000000000000000101100100111";
wait for Clk_period;

--tree 23 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011000";
Trees_din <= "00000000000000000000101110100110";
wait for Clk_period;

--tree 24 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011001";
Trees_din <= "00000000000000000000110000100101";
wait for Clk_period;

--tree 25 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011010";
Trees_din <= "00000000000000000000110010100100";
wait for Clk_period;

--tree 26 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011011";
Trees_din <= "00000000000000000000110100100011";
wait for Clk_period;

--tree 27 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011100";
Trees_din <= "00000000000000000000110110100010";
wait for Clk_period;

--tree 28 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011101";
Trees_din <= "00000000000000000000111000100001";
wait for Clk_period;

--tree 29 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011110";
Trees_din <= "00000000000000000000111010100000";
wait for Clk_period;

--tree 30 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000011111";
Trees_din <= "00000000000000000000111100011111";
wait for Clk_period;

--tree 31 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100000";
Trees_din <= "00000000000000000000111110011110";
wait for Clk_period;

--tree 32 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100001";
Trees_din <= "00000000000000000001000000011101";
wait for Clk_period;

--tree 33 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100010";
Trees_din <= "00000000000000000001000010011100";
wait for Clk_period;

--tree 34 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100011";
Trees_din <= "00000000000000000001000100011011";
wait for Clk_period;

--tree 35 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100100";
Trees_din <= "00000000000000000001000110011010";
wait for Clk_period;

--tree 36 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100101";
Trees_din <= "00000000000000000001001000011001";
wait for Clk_period;

--tree 37 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100110";
Trees_din <= "00000000000000000001001010011000";
wait for Clk_period;

--tree 38 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000100111";
Trees_din <= "00000000000000000001001100010111";
wait for Clk_period;

--tree 39 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000101000";
Trees_din <= "00000000000000000001001110010110";
wait for Clk_period;

--tree 40 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000101001";
Trees_din <= "00000000000000000001010000010101";
wait for Clk_period;

--tree 41 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000101010";
Trees_din <= "00000000000000000001010010010100";
wait for Clk_period;

--tree 42 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000101011";
Trees_din <= "00000000000000000001010100010011";
wait for Clk_period;

--tree 43 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000101100";
Trees_din <= "00000000000000000001010110010010";
wait for Clk_period;

--tree 44 belongs to class 0
-- standard deviation for this tree is 0.0
Addr <= "0000000101101";
Trees_din <= "00000000000000000001011000010001";
wait for Clk_period;

--tree 45 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000101110";
Trees_din <= "00000000000000000011011010010000";
wait for Clk_period;

--tree 46 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000101111";
Trees_din <= "00000000000000000011011100001111";
wait for Clk_period;

--tree 47 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110000";
Trees_din <= "00000000000000000011011110001110";
wait for Clk_period;

--tree 48 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110001";
Trees_din <= "00000000000000000011100000001101";
wait for Clk_period;

--tree 49 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110010";
Trees_din <= "00000000000000000011100010001100";
wait for Clk_period;

--tree 50 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110011";
Trees_din <= "00000000000000000011100100001011";
wait for Clk_period;

--tree 51 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110100";
Trees_din <= "00000000000000000011100110001010";
wait for Clk_period;

--tree 52 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110101";
Trees_din <= "00000000000000000011101000001001";
wait for Clk_period;

--tree 53 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110110";
Trees_din <= "00000000000000000011101010001000";
wait for Clk_period;

--tree 54 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000110111";
Trees_din <= "00000000000000000011101100000111";
wait for Clk_period;

--tree 55 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000111000";
Trees_din <= "00000000000000000011101110000110";
wait for Clk_period;

--tree 56 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000111001";
Trees_din <= "00000000000000000011110000000101";
wait for Clk_period;

--tree 57 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000111010";
Trees_din <= "00000000000000000011110010000100";
wait for Clk_period;

--tree 58 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000111011";
Trees_din <= "00000000000000000011110100000011";
wait for Clk_period;

--tree 59 belongs to class 1
-- standard deviation for this tree is 0.0
Addr <= "0000000111100";
Trees_din <= "00000000000000000011110110000010";
wait for Clk_period;




----------tree 0-------------------

Addr <= "0000000111101";
Trees_din <= "00000111000000000010101010000000";
wait for Clk_period;
Addr <= "0000000111110";
Trees_din <= "00000010000000000010100001000000";
wait for Clk_period;
Addr <= "0000000111111";
Trees_din <= "00000011000000000011011000100000";
wait for Clk_period;
Addr <= "0000001000000";
Trees_din <= "00000011000000000010101000010000";
wait for Clk_period;
Addr <= "0000001000001";
Trees_din <= "00000001000000000011100100001000";
wait for Clk_period;
Addr <= "0000001000010";
Trees_din <= "00000001000000000000000100000100";
wait for Clk_period;
Addr <= "0000001000011";
Trees_din <= "00000000001010000000001011110001";
wait for Clk_period;
Addr <= "0000001000100";
Trees_din <= "00000000000111010000001011110001";
wait for Clk_period;
Addr <= "0000001000101";
Trees_din <= "00000011000000000001111100000100";
wait for Clk_period;
Addr <= "0000001000110";
Trees_din <= "00000000001000000000001011110001";
wait for Clk_period;
Addr <= "0000001000111";
Trees_din <= "00000000000001110000001011110001";
wait for Clk_period;
Addr <= "0000001001000";
Trees_din <= "00000000000000000001001000001000";
wait for Clk_period;
Addr <= "0000001001001";
Trees_din <= "00000111000000000100101100000100";
wait for Clk_period;
Addr <= "0000001001010";
Trees_din <= "00000000010000110000001011110001";
wait for Clk_period;
Addr <= "0000001001011";
Trees_din <= "00000000010100110000001011110001";
wait for Clk_period;
Addr <= "0000001001100";
Trees_din <= "00000010000000000100011100000100";
wait for Clk_period;
Addr <= "0000001001101";
Trees_din <= "00000000010100010000001011110001";
wait for Clk_period;
Addr <= "0000001001110";
Trees_din <= "00000000010011100000001011110001";
wait for Clk_period;
Addr <= "0000001001111";
Trees_din <= "00000011000000000100010100010000";
wait for Clk_period;
Addr <= "0000001010000";
Trees_din <= "00000010000000000000011000001000";
wait for Clk_period;
Addr <= "0000001010001";
Trees_din <= "00000000000000000011001100000100";
wait for Clk_period;
Addr <= "0000001010010";
Trees_din <= "00000000001111010000001011110001";
wait for Clk_period;
Addr <= "0000001010011";
Trees_din <= "00000000010110100000001011110001";
wait for Clk_period;
Addr <= "0000001010100";
Trees_din <= "00000110000000000100101000000100";
wait for Clk_period;
Addr <= "0000001010101";
Trees_din <= "00000000000010000000001011110001";
wait for Clk_period;
Addr <= "0000001010110";
Trees_din <= "00000000011000000000001011110001";
wait for Clk_period;
Addr <= "0000001010111";
Trees_din <= "00000001000000000101100100001000";
wait for Clk_period;
Addr <= "0000001011000";
Trees_din <= "00000001000000000011000000000100";
wait for Clk_period;
Addr <= "0000001011001";
Trees_din <= "00000000000011000000001011110001";
wait for Clk_period;
Addr <= "0000001011010";
Trees_din <= "00000000000111010000001011110001";
wait for Clk_period;
Addr <= "0000001011011";
Trees_din <= "00000001000000000100100100000100";
wait for Clk_period;
Addr <= "0000001011100";
Trees_din <= "00000000000000000000001011110001";
wait for Clk_period;
Addr <= "0000001011101";
Trees_din <= "00000000000100010000001011110001";
wait for Clk_period;
Addr <= "0000001011110";
Trees_din <= "00000100000000000101110000100000";
wait for Clk_period;
Addr <= "0000001011111";
Trees_din <= "00000110000000000101001000010000";
wait for Clk_period;
Addr <= "0000001100000";
Trees_din <= "00000011000000000011001000001000";
wait for Clk_period;
Addr <= "0000001100001";
Trees_din <= "00000000000000000101110100000100";
wait for Clk_period;
Addr <= "0000001100010";
Trees_din <= "00000000000011010000001011110001";
wait for Clk_period;
Addr <= "0000001100011";
Trees_din <= "00000000010000010000001011110001";
wait for Clk_period;
Addr <= "0000001100100";
Trees_din <= "00000110000000000010100100000100";
wait for Clk_period;
Addr <= "0000001100101";
Trees_din <= "00000000001001110000001011110001";
wait for Clk_period;
Addr <= "0000001100110";
Trees_din <= "00000000010010000000001011110001";
wait for Clk_period;
Addr <= "0000001100111";
Trees_din <= "00000111000000000000110000001000";
wait for Clk_period;
Addr <= "0000001101000";
Trees_din <= "00000011000000000011011100000100";
wait for Clk_period;
Addr <= "0000001101001";
Trees_din <= "00000000000001110000001011110001";
wait for Clk_period;
Addr <= "0000001101010";
Trees_din <= "00000000001100010000001011110001";
wait for Clk_period;
Addr <= "0000001101011";
Trees_din <= "00000000000000000100001000000100";
wait for Clk_period;
Addr <= "0000001101100";
Trees_din <= "00000000001000110000001011110001";
wait for Clk_period;
Addr <= "0000001101101";
Trees_din <= "00000000010110000000001011110001";
wait for Clk_period;
Addr <= "0000001101110";
Trees_din <= "00000011000000000100110100010000";
wait for Clk_period;
Addr <= "0000001101111";
Trees_din <= "00000111000000000010111100001000";
wait for Clk_period;
Addr <= "0000001110000";
Trees_din <= "00000000000000000100110000000100";
wait for Clk_period;
Addr <= "0000001110001";
Trees_din <= "00000000010000110000001011110001";
wait for Clk_period;
Addr <= "0000001110010";
Trees_din <= "00000000000110100000001011110001";
wait for Clk_period;
Addr <= "0000001110011";
Trees_din <= "00000011000000000011011100000100";
wait for Clk_period;
Addr <= "0000001110100";
Trees_din <= "00000000010000000000001011110001";
wait for Clk_period;
Addr <= "0000001110101";
Trees_din <= "00000000001110100000001011110001";
wait for Clk_period;
Addr <= "0000001110110";
Trees_din <= "00000100000000000001000000001000";
wait for Clk_period;
Addr <= "0000001110111";
Trees_din <= "00000101000000000100001100000100";
wait for Clk_period;
Addr <= "0000001111000";
Trees_din <= "00000000010000100000001011110001";
wait for Clk_period;
Addr <= "0000001111001";
Trees_din <= "00000000000111100000001011110001";
wait for Clk_period;
Addr <= "0000001111010";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "0000001111011";
Trees_din <= "00000000010110010000001011110001";
wait for Clk_period;
Addr <= "0000001111100";
Trees_din <= "00000000000101010000001011110001";
wait for Clk_period;
Addr <= "0000001111101";
Trees_din <= "00000100000000000100011001000000";
wait for Clk_period;
Addr <= "0000001111110";
Trees_din <= "00000111000000000101101100100000";
wait for Clk_period;
Addr <= "0000001111111";
Trees_din <= "00000111000000000100111100010000";
wait for Clk_period;
Addr <= "0000010000000";
Trees_din <= "00000010000000000000110100001000";
wait for Clk_period;
Addr <= "0000010000001";
Trees_din <= "00000000000000000000101000000100";
wait for Clk_period;
Addr <= "0000010000010";
Trees_din <= "00000000000110010000001011110001";
wait for Clk_period;
Addr <= "0000010000011";
Trees_din <= "00000000000110000000001011110001";
wait for Clk_period;
Addr <= "0000010000100";
Trees_din <= "00000001000000000010100000000100";
wait for Clk_period;
Addr <= "0000010000101";
Trees_din <= "00000000000110100000001011110001";
wait for Clk_period;
Addr <= "0000010000110";
Trees_din <= "00000000000010000000001011110001";
wait for Clk_period;
Addr <= "0000010000111";
Trees_din <= "00000001000000000000011100001000";
wait for Clk_period;
Addr <= "0000010001000";
Trees_din <= "00000100000000000101001000000100";
wait for Clk_period;
Addr <= "0000010001001";
Trees_din <= "00000000010101110000001011110001";
wait for Clk_period;
Addr <= "0000010001010";
Trees_din <= "00000000000001010000001011110001";
wait for Clk_period;
Addr <= "0000010001011";
Trees_din <= "00000000000000000110001100000100";
wait for Clk_period;
Addr <= "0000010001100";
Trees_din <= "00000000010011110000001011110001";
wait for Clk_period;
Addr <= "0000010001101";
Trees_din <= "00000000001001100000001011110001";
wait for Clk_period;
Addr <= "0000010001110";
Trees_din <= "00000110000000000100110100010000";
wait for Clk_period;
Addr <= "0000010001111";
Trees_din <= "00000110000000000110001000001000";
wait for Clk_period;
Addr <= "0000010010000";
Trees_din <= "00000101000000000000111000000100";
wait for Clk_period;
Addr <= "0000010010001";
Trees_din <= "00000000000000010000001011110001";
wait for Clk_period;
Addr <= "0000010010010";
Trees_din <= "00000000010100100000001011110001";
wait for Clk_period;
Addr <= "0000010010011";
Trees_din <= "00000010000000000110000100000100";
wait for Clk_period;
Addr <= "0000010010100";
Trees_din <= "00000000001010000000001011110001";
wait for Clk_period;
Addr <= "0000010010101";
Trees_din <= "00000000000101100000001011110001";
wait for Clk_period;
Addr <= "0000010010110";
Trees_din <= "00000100000000000000001100001000";
wait for Clk_period;
Addr <= "0000010010111";
Trees_din <= "00000100000000000001100000000100";
wait for Clk_period;
Addr <= "0000010011000";
Trees_din <= "00000000000011010000001011110001";
wait for Clk_period;
Addr <= "0000010011001";
Trees_din <= "00000000010001110000001011110001";
wait for Clk_period;
Addr <= "0000010011010";
Trees_din <= "00000111000000000010110100000100";
wait for Clk_period;
Addr <= "0000010011011";
Trees_din <= "00000000001010000000001011110001";
wait for Clk_period;
Addr <= "0000010011100";
Trees_din <= "00000000000001100000001011110001";
wait for Clk_period;
Addr <= "0000010011101";
Trees_din <= "00000000000000000100101100100000";
wait for Clk_period;
Addr <= "0000010011110";
Trees_din <= "00000010000000000110010000010000";
wait for Clk_period;
Addr <= "0000010011111";
Trees_din <= "00000111000000000001000000001000";
wait for Clk_period;
Addr <= "0000010100000";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "0000010100001";
Trees_din <= "00000000001101110000001011110001";
wait for Clk_period;
Addr <= "0000010100010";
Trees_din <= "00000000000101000000001011110001";
wait for Clk_period;
Addr <= "0000010100011";
Trees_din <= "00000001000000000100101000000100";
wait for Clk_period;
Addr <= "0000010100100";
Trees_din <= "00000000000111000000001011110001";
wait for Clk_period;
Addr <= "0000010100101";
Trees_din <= "00000000001100000000001011110001";
wait for Clk_period;
Addr <= "0000010100110";
Trees_din <= "00000000000000000001011000001000";
wait for Clk_period;
Addr <= "0000010100111";
Trees_din <= "00000000000000000110010000000100";
wait for Clk_period;
Addr <= "0000010101000";
Trees_din <= "00000000010001010000001011110001";
wait for Clk_period;
Addr <= "0000010101001";
Trees_din <= "00000000010000000000001011110001";
wait for Clk_period;
Addr <= "0000010101010";
Trees_din <= "00000101000000000011100000000100";
wait for Clk_period;
Addr <= "0000010101011";
Trees_din <= "00000000000101100000001011110001";
wait for Clk_period;
Addr <= "0000010101100";
Trees_din <= "00000000010100010000001011110001";
wait for Clk_period;
Addr <= "0000010101101";
Trees_din <= "00000011000000000011100000010000";
wait for Clk_period;
Addr <= "0000010101110";
Trees_din <= "00000101000000000100000000001000";
wait for Clk_period;
Addr <= "0000010101111";
Trees_din <= "00000111000000000011100000000100";
wait for Clk_period;
Addr <= "0000010110000";
Trees_din <= "00000000001100100000001011110001";
wait for Clk_period;
Addr <= "0000010110001";
Trees_din <= "00000000010011100000001011110001";
wait for Clk_period;
Addr <= "0000010110010";
Trees_din <= "00000110000000000001010100000100";
wait for Clk_period;
Addr <= "0000010110011";
Trees_din <= "00000000000111100000001011110001";
wait for Clk_period;
Addr <= "0000010110100";
Trees_din <= "00000000001001000000001011110001";
wait for Clk_period;
Addr <= "0000010110101";
Trees_din <= "00000010000000000101100100001000";
wait for Clk_period;
Addr <= "0000010110110";
Trees_din <= "00000111000000000010010000000100";
wait for Clk_period;
Addr <= "0000010110111";
Trees_din <= "00000000000111100000001011110001";
wait for Clk_period;
Addr <= "0000010111000";
Trees_din <= "00000000010111100000001011110001";
wait for Clk_period;
Addr <= "0000010111001";
Trees_din <= "00000101000000000000000000000100";
wait for Clk_period;
Addr <= "0000010111010";
Trees_din <= "00000000010110010000001011110001";
wait for Clk_period;
Addr <= "0000010111011";
Trees_din <= "00000000000001000000001011110001";
wait for Clk_period;



----------tree 1-------------------

Addr <= "0000010111100";
Trees_din <= "00000111000000000100110110000000";
wait for Clk_period;
Addr <= "0000010111101";
Trees_din <= "00000100000000000100011101000000";
wait for Clk_period;
Addr <= "0000010111110";
Trees_din <= "00000000000000000011010100100000";
wait for Clk_period;
Addr <= "0000010111111";
Trees_din <= "00000111000000000011111000010000";
wait for Clk_period;
Addr <= "0000011000000";
Trees_din <= "00000010000000000011000100001000";
wait for Clk_period;
Addr <= "0000011000001";
Trees_din <= "00000111000000000000001000000100";
wait for Clk_period;
Addr <= "0000011000010";
Trees_din <= "00000000000111100000010011101101";
wait for Clk_period;
Addr <= "0000011000011";
Trees_din <= "00000000001110010000010011101101";
wait for Clk_period;
Addr <= "0000011000100";
Trees_din <= "00000101000000000100110100000100";
wait for Clk_period;
Addr <= "0000011000101";
Trees_din <= "00000000010100110000010011101101";
wait for Clk_period;
Addr <= "0000011000110";
Trees_din <= "00000000000011100000010011101101";
wait for Clk_period;
Addr <= "0000011000111";
Trees_din <= "00000100000000000011010000001000";
wait for Clk_period;
Addr <= "0000011001000";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "0000011001001";
Trees_din <= "00000000001001110000010011101101";
wait for Clk_period;
Addr <= "0000011001010";
Trees_din <= "00000000010000100000010011101101";
wait for Clk_period;
Addr <= "0000011001011";
Trees_din <= "00000100000000000010011100000100";
wait for Clk_period;
Addr <= "0000011001100";
Trees_din <= "00000000001111110000010011101101";
wait for Clk_period;
Addr <= "0000011001101";
Trees_din <= "00000000010101010000010011101101";
wait for Clk_period;
Addr <= "0000011001110";
Trees_din <= "00000101000000000000101100010000";
wait for Clk_period;
Addr <= "0000011001111";
Trees_din <= "00000110000000000000110000001000";
wait for Clk_period;
Addr <= "0000011010000";
Trees_din <= "00000010000000000000111100000100";
wait for Clk_period;
Addr <= "0000011010001";
Trees_din <= "00000000001101000000010011101101";
wait for Clk_period;
Addr <= "0000011010010";
Trees_din <= "00000000000100110000010011101101";
wait for Clk_period;
Addr <= "0000011010011";
Trees_din <= "00000110000000000001011100000100";
wait for Clk_period;
Addr <= "0000011010100";
Trees_din <= "00000000010100010000010011101101";
wait for Clk_period;
Addr <= "0000011010101";
Trees_din <= "00000000000111110000010011101101";
wait for Clk_period;
Addr <= "0000011010110";
Trees_din <= "00000111000000000101010100001000";
wait for Clk_period;
Addr <= "0000011010111";
Trees_din <= "00000010000000000010111100000100";
wait for Clk_period;
Addr <= "0000011011000";
Trees_din <= "00000000001101100000010011101101";
wait for Clk_period;
Addr <= "0000011011001";
Trees_din <= "00000000001001000000010011101101";
wait for Clk_period;
Addr <= "0000011011010";
Trees_din <= "00000011000000000110000100000100";
wait for Clk_period;
Addr <= "0000011011011";
Trees_din <= "00000000010110100000010011101101";
wait for Clk_period;
Addr <= "0000011011100";
Trees_din <= "00000000000010100000010011101101";
wait for Clk_period;
Addr <= "0000011011101";
Trees_din <= "00000100000000000000011100100000";
wait for Clk_period;
Addr <= "0000011011110";
Trees_din <= "00000010000000000011111000010000";
wait for Clk_period;
Addr <= "0000011011111";
Trees_din <= "00000101000000000100101100001000";
wait for Clk_period;
Addr <= "0000011100000";
Trees_din <= "00000110000000000110001000000100";
wait for Clk_period;
Addr <= "0000011100001";
Trees_din <= "00000000001100110000010011101101";
wait for Clk_period;
Addr <= "0000011100010";
Trees_din <= "00000000010001100000010011101101";
wait for Clk_period;
Addr <= "0000011100011";
Trees_din <= "00000001000000000010100100000100";
wait for Clk_period;
Addr <= "0000011100100";
Trees_din <= "00000000001101000000010011101101";
wait for Clk_period;
Addr <= "0000011100101";
Trees_din <= "00000000001110100000010011101101";
wait for Clk_period;
Addr <= "0000011100110";
Trees_din <= "00000011000000000101001100001000";
wait for Clk_period;
Addr <= "0000011100111";
Trees_din <= "00000010000000000010001100000100";
wait for Clk_period;
Addr <= "0000011101000";
Trees_din <= "00000000000011000000010011101101";
wait for Clk_period;
Addr <= "0000011101001";
Trees_din <= "00000000001001000000010011101101";
wait for Clk_period;
Addr <= "0000011101010";
Trees_din <= "00000111000000000010110000000100";
wait for Clk_period;
Addr <= "0000011101011";
Trees_din <= "00000000000001010000010011101101";
wait for Clk_period;
Addr <= "0000011101100";
Trees_din <= "00000000001001010000010011101101";
wait for Clk_period;
Addr <= "0000011101101";
Trees_din <= "00000110000000000010101100010000";
wait for Clk_period;
Addr <= "0000011101110";
Trees_din <= "00000100000000000000011100001000";
wait for Clk_period;
Addr <= "0000011101111";
Trees_din <= "00000110000000000101011000000100";
wait for Clk_period;
Addr <= "0000011110000";
Trees_din <= "00000000011000000000010011101101";
wait for Clk_period;
Addr <= "0000011110001";
Trees_din <= "00000000000100110000010011101101";
wait for Clk_period;
Addr <= "0000011110010";
Trees_din <= "00000010000000000010011100000100";
wait for Clk_period;
Addr <= "0000011110011";
Trees_din <= "00000000011000110000010011101101";
wait for Clk_period;
Addr <= "0000011110100";
Trees_din <= "00000000010100100000010011101101";
wait for Clk_period;
Addr <= "0000011110101";
Trees_din <= "00000001000000000001110100001000";
wait for Clk_period;
Addr <= "0000011110110";
Trees_din <= "00000100000000000000101100000100";
wait for Clk_period;
Addr <= "0000011110111";
Trees_din <= "00000000001111000000010011101101";
wait for Clk_period;
Addr <= "0000011111000";
Trees_din <= "00000000001011010000010011101101";
wait for Clk_period;
Addr <= "0000011111001";
Trees_din <= "00000111000000000001111100000100";
wait for Clk_period;
Addr <= "0000011111010";
Trees_din <= "00000000010001010000010011101101";
wait for Clk_period;
Addr <= "0000011111011";
Trees_din <= "00000000010101100000010011101101";
wait for Clk_period;
Addr <= "0000011111100";
Trees_din <= "00000000000000000001000101000000";
wait for Clk_period;
Addr <= "0000011111101";
Trees_din <= "00000101000000000001000000100000";
wait for Clk_period;
Addr <= "0000011111110";
Trees_din <= "00000010000000000001010100010000";
wait for Clk_period;
Addr <= "0000011111111";
Trees_din <= "00000011000000000000111000001000";
wait for Clk_period;
Addr <= "0000100000000";
Trees_din <= "00000010000000000001111000000100";
wait for Clk_period;
Addr <= "0000100000001";
Trees_din <= "00000000010110000000010011101101";
wait for Clk_period;
Addr <= "0000100000010";
Trees_din <= "00000000010101100000010011101101";
wait for Clk_period;
Addr <= "0000100000011";
Trees_din <= "00000101000000000011011100000100";
wait for Clk_period;
Addr <= "0000100000100";
Trees_din <= "00000000001000110000010011101101";
wait for Clk_period;
Addr <= "0000100000101";
Trees_din <= "00000000010011100000010011101101";
wait for Clk_period;
Addr <= "0000100000110";
Trees_din <= "00000110000000000000001100001000";
wait for Clk_period;
Addr <= "0000100000111";
Trees_din <= "00000001000000000101101000000100";
wait for Clk_period;
Addr <= "0000100001000";
Trees_din <= "00000000001011010000010011101101";
wait for Clk_period;
Addr <= "0000100001001";
Trees_din <= "00000000011000010000010011101101";
wait for Clk_period;
Addr <= "0000100001010";
Trees_din <= "00000101000000000100111000000100";
wait for Clk_period;
Addr <= "0000100001011";
Trees_din <= "00000000001011100000010011101101";
wait for Clk_period;
Addr <= "0000100001100";
Trees_din <= "00000000000010010000010011101101";
wait for Clk_period;
Addr <= "0000100001101";
Trees_din <= "00000101000000000110000100010000";
wait for Clk_period;
Addr <= "0000100001110";
Trees_din <= "00000110000000000000110000001000";
wait for Clk_period;
Addr <= "0000100001111";
Trees_din <= "00000001000000000000011000000100";
wait for Clk_period;
Addr <= "0000100010000";
Trees_din <= "00000000000010110000010011101101";
wait for Clk_period;
Addr <= "0000100010001";
Trees_din <= "00000000011001000000010011101101";
wait for Clk_period;
Addr <= "0000100010010";
Trees_din <= "00000100000000000011011100000100";
wait for Clk_period;
Addr <= "0000100010011";
Trees_din <= "00000000010000000000010011101101";
wait for Clk_period;
Addr <= "0000100010100";
Trees_din <= "00000000000010010000010011101101";
wait for Clk_period;
Addr <= "0000100010101";
Trees_din <= "00000101000000000110001000001000";
wait for Clk_period;
Addr <= "0000100010110";
Trees_din <= "00000100000000000101001100000100";
wait for Clk_period;
Addr <= "0000100010111";
Trees_din <= "00000000010101000000010011101101";
wait for Clk_period;
Addr <= "0000100011000";
Trees_din <= "00000000010001010000010011101101";
wait for Clk_period;
Addr <= "0000100011001";
Trees_din <= "00000000000000000001000100000100";
wait for Clk_period;
Addr <= "0000100011010";
Trees_din <= "00000000001011010000010011101101";
wait for Clk_period;
Addr <= "0000100011011";
Trees_din <= "00000000001101010000010011101101";
wait for Clk_period;
Addr <= "0000100011100";
Trees_din <= "00000111000000000010000000100000";
wait for Clk_period;
Addr <= "0000100011101";
Trees_din <= "00000101000000000100100000010000";
wait for Clk_period;
Addr <= "0000100011110";
Trees_din <= "00000111000000000001001100001000";
wait for Clk_period;
Addr <= "0000100011111";
Trees_din <= "00000101000000000011110100000100";
wait for Clk_period;
Addr <= "0000100100000";
Trees_din <= "00000000001011110000010011101101";
wait for Clk_period;
Addr <= "0000100100001";
Trees_din <= "00000000001101000000010011101101";
wait for Clk_period;
Addr <= "0000100100010";
Trees_din <= "00000010000000000100001100000100";
wait for Clk_period;
Addr <= "0000100100011";
Trees_din <= "00000000001000110000010011101101";
wait for Clk_period;
Addr <= "0000100100100";
Trees_din <= "00000000001010000000010011101101";
wait for Clk_period;
Addr <= "0000100100101";
Trees_din <= "00000011000000000001110000001000";
wait for Clk_period;
Addr <= "0000100100110";
Trees_din <= "00000110000000000101000000000100";
wait for Clk_period;
Addr <= "0000100100111";
Trees_din <= "00000000010011110000010011101101";
wait for Clk_period;
Addr <= "0000100101000";
Trees_din <= "00000000001100010000010011101101";
wait for Clk_period;
Addr <= "0000100101001";
Trees_din <= "00000101000000000100110100000100";
wait for Clk_period;
Addr <= "0000100101010";
Trees_din <= "00000000010100100000010011101101";
wait for Clk_period;
Addr <= "0000100101011";
Trees_din <= "00000000000011110000010011101101";
wait for Clk_period;
Addr <= "0000100101100";
Trees_din <= "00000101000000000011110000010000";
wait for Clk_period;
Addr <= "0000100101101";
Trees_din <= "00000011000000000001011000001000";
wait for Clk_period;
Addr <= "0000100101110";
Trees_din <= "00000100000000000011011000000100";
wait for Clk_period;
Addr <= "0000100101111";
Trees_din <= "00000000001100100000010011101101";
wait for Clk_period;
Addr <= "0000100110000";
Trees_din <= "00000000001001010000010011101101";
wait for Clk_period;
Addr <= "0000100110001";
Trees_din <= "00000111000000000100001000000100";
wait for Clk_period;
Addr <= "0000100110010";
Trees_din <= "00000000010110010000010011101101";
wait for Clk_period;
Addr <= "0000100110011";
Trees_din <= "00000000010000000000010011101101";
wait for Clk_period;
Addr <= "0000100110100";
Trees_din <= "00000011000000000100111000001000";
wait for Clk_period;
Addr <= "0000100110101";
Trees_din <= "00000011000000000000000000000100";
wait for Clk_period;
Addr <= "0000100110110";
Trees_din <= "00000000000011110000010011101101";
wait for Clk_period;
Addr <= "0000100110111";
Trees_din <= "00000000011001000000010011101101";
wait for Clk_period;
Addr <= "0000100111000";
Trees_din <= "00000101000000000100100100000100";
wait for Clk_period;
Addr <= "0000100111001";
Trees_din <= "00000000001011100000010011101101";
wait for Clk_period;
Addr <= "0000100111010";
Trees_din <= "00000000010011110000010011101101";
wait for Clk_period;



----------tree 2-------------------

Addr <= "0000100111011";
Trees_din <= "00000100000000000000111010000000";
wait for Clk_period;
Addr <= "0000100111100";
Trees_din <= "00000110000000000100110101000000";
wait for Clk_period;
Addr <= "0000100111101";
Trees_din <= "00000001000000000010110100100000";
wait for Clk_period;
Addr <= "0000100111110";
Trees_din <= "00000101000000000101001000010000";
wait for Clk_period;
Addr <= "0000100111111";
Trees_din <= "00000010000000000010110000001000";
wait for Clk_period;
Addr <= "0000101000000";
Trees_din <= "00000010000000000100001100000100";
wait for Clk_period;
Addr <= "0000101000001";
Trees_din <= "00000000000011100000011011101001";
wait for Clk_period;
Addr <= "0000101000010";
Trees_din <= "00000000010011000000011011101001";
wait for Clk_period;
Addr <= "0000101000011";
Trees_din <= "00000111000000000011000100000100";
wait for Clk_period;
Addr <= "0000101000100";
Trees_din <= "00000000010001100000011011101001";
wait for Clk_period;
Addr <= "0000101000101";
Trees_din <= "00000000001000100000011011101001";
wait for Clk_period;
Addr <= "0000101000110";
Trees_din <= "00000101000000000001100000001000";
wait for Clk_period;
Addr <= "0000101000111";
Trees_din <= "00000010000000000100011000000100";
wait for Clk_period;
Addr <= "0000101001000";
Trees_din <= "00000000010111110000011011101001";
wait for Clk_period;
Addr <= "0000101001001";
Trees_din <= "00000000001000000000011011101001";
wait for Clk_period;
Addr <= "0000101001010";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "0000101001011";
Trees_din <= "00000000010010000000011011101001";
wait for Clk_period;
Addr <= "0000101001100";
Trees_din <= "00000000010100110000011011101001";
wait for Clk_period;
Addr <= "0000101001101";
Trees_din <= "00000011000000000010111000010000";
wait for Clk_period;
Addr <= "0000101001110";
Trees_din <= "00000010000000000101100100001000";
wait for Clk_period;
Addr <= "0000101001111";
Trees_din <= "00000000000000000011001000000100";
wait for Clk_period;
Addr <= "0000101010000";
Trees_din <= "00000000001111100000011011101001";
wait for Clk_period;
Addr <= "0000101010001";
Trees_din <= "00000000000001000000011011101001";
wait for Clk_period;
Addr <= "0000101010010";
Trees_din <= "00000000000000000011110100000100";
wait for Clk_period;
Addr <= "0000101010011";
Trees_din <= "00000000010010100000011011101001";
wait for Clk_period;
Addr <= "0000101010100";
Trees_din <= "00000000000011110000011011101001";
wait for Clk_period;
Addr <= "0000101010101";
Trees_din <= "00000001000000000100010000001000";
wait for Clk_period;
Addr <= "0000101010110";
Trees_din <= "00000101000000000001110000000100";
wait for Clk_period;
Addr <= "0000101010111";
Trees_din <= "00000000001000110000011011101001";
wait for Clk_period;
Addr <= "0000101011000";
Trees_din <= "00000000000001110000011011101001";
wait for Clk_period;
Addr <= "0000101011001";
Trees_din <= "00000000000000000001000000000100";
wait for Clk_period;
Addr <= "0000101011010";
Trees_din <= "00000000001011000000011011101001";
wait for Clk_period;
Addr <= "0000101011011";
Trees_din <= "00000000010111000000011011101001";
wait for Clk_period;
Addr <= "0000101011100";
Trees_din <= "00000001000000000100001100100000";
wait for Clk_period;
Addr <= "0000101011101";
Trees_din <= "00000101000000000001000100010000";
wait for Clk_period;
Addr <= "0000101011110";
Trees_din <= "00000010000000000101100100001000";
wait for Clk_period;
Addr <= "0000101011111";
Trees_din <= "00000000000000000001001000000100";
wait for Clk_period;
Addr <= "0000101100000";
Trees_din <= "00000000011000100000011011101001";
wait for Clk_period;
Addr <= "0000101100001";
Trees_din <= "00000000010101110000011011101001";
wait for Clk_period;
Addr <= "0000101100010";
Trees_din <= "00000010000000000000111100000100";
wait for Clk_period;
Addr <= "0000101100011";
Trees_din <= "00000000011000010000011011101001";
wait for Clk_period;
Addr <= "0000101100100";
Trees_din <= "00000000010011100000011011101001";
wait for Clk_period;
Addr <= "0000101100101";
Trees_din <= "00000110000000000010010000001000";
wait for Clk_period;
Addr <= "0000101100110";
Trees_din <= "00000011000000000011110100000100";
wait for Clk_period;
Addr <= "0000101100111";
Trees_din <= "00000000010110100000011011101001";
wait for Clk_period;
Addr <= "0000101101000";
Trees_din <= "00000000001111010000011011101001";
wait for Clk_period;
Addr <= "0000101101001";
Trees_din <= "00000011000000000110010000000100";
wait for Clk_period;
Addr <= "0000101101010";
Trees_din <= "00000000000110110000011011101001";
wait for Clk_period;
Addr <= "0000101101011";
Trees_din <= "00000000010101000000011011101001";
wait for Clk_period;
Addr <= "0000101101100";
Trees_din <= "00000110000000000101011100010000";
wait for Clk_period;
Addr <= "0000101101101";
Trees_din <= "00000001000000000000110000001000";
wait for Clk_period;
Addr <= "0000101101110";
Trees_din <= "00000110000000000000100100000100";
wait for Clk_period;
Addr <= "0000101101111";
Trees_din <= "00000000001101110000011011101001";
wait for Clk_period;
Addr <= "0000101110000";
Trees_din <= "00000000000100010000011011101001";
wait for Clk_period;
Addr <= "0000101110001";
Trees_din <= "00000111000000000101111100000100";
wait for Clk_period;
Addr <= "0000101110010";
Trees_din <= "00000000001100100000011011101001";
wait for Clk_period;
Addr <= "0000101110011";
Trees_din <= "00000000010001100000011011101001";
wait for Clk_period;
Addr <= "0000101110100";
Trees_din <= "00000011000000000100001000001000";
wait for Clk_period;
Addr <= "0000101110101";
Trees_din <= "00000100000000000101011000000100";
wait for Clk_period;
Addr <= "0000101110110";
Trees_din <= "00000000000010010000011011101001";
wait for Clk_period;
Addr <= "0000101110111";
Trees_din <= "00000000000110000000011011101001";
wait for Clk_period;
Addr <= "0000101111000";
Trees_din <= "00000110000000000010111000000100";
wait for Clk_period;
Addr <= "0000101111001";
Trees_din <= "00000000000000110000011011101001";
wait for Clk_period;
Addr <= "0000101111010";
Trees_din <= "00000000010010000000011011101001";
wait for Clk_period;
Addr <= "0000101111011";
Trees_din <= "00000000000000000010101101000000";
wait for Clk_period;
Addr <= "0000101111100";
Trees_din <= "00000000000000000000111100100000";
wait for Clk_period;
Addr <= "0000101111101";
Trees_din <= "00000111000000000001111100010000";
wait for Clk_period;
Addr <= "0000101111110";
Trees_din <= "00000110000000000010000000001000";
wait for Clk_period;
Addr <= "0000101111111";
Trees_din <= "00000100000000000001100000000100";
wait for Clk_period;
Addr <= "0000110000000";
Trees_din <= "00000000011000010000011011101001";
wait for Clk_period;
Addr <= "0000110000001";
Trees_din <= "00000000000101100000011011101001";
wait for Clk_period;
Addr <= "0000110000010";
Trees_din <= "00000000000000000001010000000100";
wait for Clk_period;
Addr <= "0000110000011";
Trees_din <= "00000000010011000000011011101001";
wait for Clk_period;
Addr <= "0000110000100";
Trees_din <= "00000000001101110000011011101001";
wait for Clk_period;
Addr <= "0000110000101";
Trees_din <= "00000011000000000100110000001000";
wait for Clk_period;
Addr <= "0000110000110";
Trees_din <= "00000011000000000101001000000100";
wait for Clk_period;
Addr <= "0000110000111";
Trees_din <= "00000000001100010000011011101001";
wait for Clk_period;
Addr <= "0000110001000";
Trees_din <= "00000000000111100000011011101001";
wait for Clk_period;
Addr <= "0000110001001";
Trees_din <= "00000010000000000010100000000100";
wait for Clk_period;
Addr <= "0000110001010";
Trees_din <= "00000000010010000000011011101001";
wait for Clk_period;
Addr <= "0000110001011";
Trees_din <= "00000000000001110000011011101001";
wait for Clk_period;
Addr <= "0000110001100";
Trees_din <= "00000000000000000010101000010000";
wait for Clk_period;
Addr <= "0000110001101";
Trees_din <= "00000011000000000001111000001000";
wait for Clk_period;
Addr <= "0000110001110";
Trees_din <= "00000111000000000100110000000100";
wait for Clk_period;
Addr <= "0000110001111";
Trees_din <= "00000000000011110000011011101001";
wait for Clk_period;
Addr <= "0000110010000";
Trees_din <= "00000000010011110000011011101001";
wait for Clk_period;
Addr <= "0000110010001";
Trees_din <= "00000011000000000101001100000100";
wait for Clk_period;
Addr <= "0000110010010";
Trees_din <= "00000000000111110000011011101001";
wait for Clk_period;
Addr <= "0000110010011";
Trees_din <= "00000000000001010000011011101001";
wait for Clk_period;
Addr <= "0000110010100";
Trees_din <= "00000100000000000101100000001000";
wait for Clk_period;
Addr <= "0000110010101";
Trees_din <= "00000111000000000010101000000100";
wait for Clk_period;
Addr <= "0000110010110";
Trees_din <= "00000000001011000000011011101001";
wait for Clk_period;
Addr <= "0000110010111";
Trees_din <= "00000000001101100000011011101001";
wait for Clk_period;
Addr <= "0000110011000";
Trees_din <= "00000001000000000000001000000100";
wait for Clk_period;
Addr <= "0000110011001";
Trees_din <= "00000000000110100000011011101001";
wait for Clk_period;
Addr <= "0000110011010";
Trees_din <= "00000000000000100000011011101001";
wait for Clk_period;
Addr <= "0000110011011";
Trees_din <= "00000101000000000101110000100000";
wait for Clk_period;
Addr <= "0000110011100";
Trees_din <= "00000011000000000101011100010000";
wait for Clk_period;
Addr <= "0000110011101";
Trees_din <= "00000111000000000101110000001000";
wait for Clk_period;
Addr <= "0000110011110";
Trees_din <= "00000001000000000011110000000100";
wait for Clk_period;
Addr <= "0000110011111";
Trees_din <= "00000000001110110000011011101001";
wait for Clk_period;
Addr <= "0000110100000";
Trees_din <= "00000000010101110000011011101001";
wait for Clk_period;
Addr <= "0000110100001";
Trees_din <= "00000000000000000110001100000100";
wait for Clk_period;
Addr <= "0000110100010";
Trees_din <= "00000000010010000000011011101001";
wait for Clk_period;
Addr <= "0000110100011";
Trees_din <= "00000000010101010000011011101001";
wait for Clk_period;
Addr <= "0000110100100";
Trees_din <= "00000000000000000001000100001000";
wait for Clk_period;
Addr <= "0000110100101";
Trees_din <= "00000101000000000000101000000100";
wait for Clk_period;
Addr <= "0000110100110";
Trees_din <= "00000000001101000000011011101001";
wait for Clk_period;
Addr <= "0000110100111";
Trees_din <= "00000000000010010000011011101001";
wait for Clk_period;
Addr <= "0000110101000";
Trees_din <= "00000001000000000100010000000100";
wait for Clk_period;
Addr <= "0000110101001";
Trees_din <= "00000000011000100000011011101001";
wait for Clk_period;
Addr <= "0000110101010";
Trees_din <= "00000000001000000000011011101001";
wait for Clk_period;
Addr <= "0000110101011";
Trees_din <= "00000100000000000001100100010000";
wait for Clk_period;
Addr <= "0000110101100";
Trees_din <= "00000010000000000101001000001000";
wait for Clk_period;
Addr <= "0000110101101";
Trees_din <= "00000110000000000000110000000100";
wait for Clk_period;
Addr <= "0000110101110";
Trees_din <= "00000000001010110000011011101001";
wait for Clk_period;
Addr <= "0000110101111";
Trees_din <= "00000000001001010000011011101001";
wait for Clk_period;
Addr <= "0000110110000";
Trees_din <= "00000000000000000011001100000100";
wait for Clk_period;
Addr <= "0000110110001";
Trees_din <= "00000000000111100000011011101001";
wait for Clk_period;
Addr <= "0000110110010";
Trees_din <= "00000000000011100000011011101001";
wait for Clk_period;
Addr <= "0000110110011";
Trees_din <= "00000110000000000011101100001000";
wait for Clk_period;
Addr <= "0000110110100";
Trees_din <= "00000110000000000000001000000100";
wait for Clk_period;
Addr <= "0000110110101";
Trees_din <= "00000000000001010000011011101001";
wait for Clk_period;
Addr <= "0000110110110";
Trees_din <= "00000000001101000000011011101001";
wait for Clk_period;
Addr <= "0000110110111";
Trees_din <= "00000011000000000100110100000100";
wait for Clk_period;
Addr <= "0000110111000";
Trees_din <= "00000000000101100000011011101001";
wait for Clk_period;
Addr <= "0000110111001";
Trees_din <= "00000000010110010000011011101001";
wait for Clk_period;



----------tree 3-------------------

Addr <= "0000110111010";
Trees_din <= "00000111000000000001010110000000";
wait for Clk_period;
Addr <= "0000110111011";
Trees_din <= "00000001000000000011101001000000";
wait for Clk_period;
Addr <= "0000110111100";
Trees_din <= "00000111000000000101001100100000";
wait for Clk_period;
Addr <= "0000110111101";
Trees_din <= "00000000000000000010110000010000";
wait for Clk_period;
Addr <= "0000110111110";
Trees_din <= "00000110000000000101110000001000";
wait for Clk_period;
Addr <= "0000110111111";
Trees_din <= "00000001000000000000100100000100";
wait for Clk_period;
Addr <= "0000111000000";
Trees_din <= "00000000010101100000100011100101";
wait for Clk_period;
Addr <= "0000111000001";
Trees_din <= "00000000001011110000100011100101";
wait for Clk_period;
Addr <= "0000111000010";
Trees_din <= "00000001000000000010010100000100";
wait for Clk_period;
Addr <= "0000111000011";
Trees_din <= "00000000001110110000100011100101";
wait for Clk_period;
Addr <= "0000111000100";
Trees_din <= "00000000001000110000100011100101";
wait for Clk_period;
Addr <= "0000111000101";
Trees_din <= "00000010000000000100101100001000";
wait for Clk_period;
Addr <= "0000111000110";
Trees_din <= "00000000000000000011011000000100";
wait for Clk_period;
Addr <= "0000111000111";
Trees_din <= "00000000000001110000100011100101";
wait for Clk_period;
Addr <= "0000111001000";
Trees_din <= "00000000001011110000100011100101";
wait for Clk_period;
Addr <= "0000111001001";
Trees_din <= "00000000000000000101101100000100";
wait for Clk_period;
Addr <= "0000111001010";
Trees_din <= "00000000010100010000100011100101";
wait for Clk_period;
Addr <= "0000111001011";
Trees_din <= "00000000010100110000100011100101";
wait for Clk_period;
Addr <= "0000111001100";
Trees_din <= "00000100000000000000101100010000";
wait for Clk_period;
Addr <= "0000111001101";
Trees_din <= "00000111000000000000101000001000";
wait for Clk_period;
Addr <= "0000111001110";
Trees_din <= "00000000000000000110000100000100";
wait for Clk_period;
Addr <= "0000111001111";
Trees_din <= "00000000010110110000100011100101";
wait for Clk_period;
Addr <= "0000111010000";
Trees_din <= "00000000001000110000100011100101";
wait for Clk_period;
Addr <= "0000111010001";
Trees_din <= "00000100000000000110000000000100";
wait for Clk_period;
Addr <= "0000111010010";
Trees_din <= "00000000000110010000100011100101";
wait for Clk_period;
Addr <= "0000111010011";
Trees_din <= "00000000010000010000100011100101";
wait for Clk_period;
Addr <= "0000111010100";
Trees_din <= "00000001000000000100100100001000";
wait for Clk_period;
Addr <= "0000111010101";
Trees_din <= "00000011000000000010010100000100";
wait for Clk_period;
Addr <= "0000111010110";
Trees_din <= "00000000001011010000100011100101";
wait for Clk_period;
Addr <= "0000111010111";
Trees_din <= "00000000000110000000100011100101";
wait for Clk_period;
Addr <= "0000111011000";
Trees_din <= "00000010000000000101101000000100";
wait for Clk_period;
Addr <= "0000111011001";
Trees_din <= "00000000000011110000100011100101";
wait for Clk_period;
Addr <= "0000111011010";
Trees_din <= "00000000010001100000100011100101";
wait for Clk_period;
Addr <= "0000111011011";
Trees_din <= "00000011000000000010011000100000";
wait for Clk_period;
Addr <= "0000111011100";
Trees_din <= "00000111000000000000100000010000";
wait for Clk_period;
Addr <= "0000111011101";
Trees_din <= "00000010000000000101010000001000";
wait for Clk_period;
Addr <= "0000111011110";
Trees_din <= "00000101000000000001001100000100";
wait for Clk_period;
Addr <= "0000111011111";
Trees_din <= "00000000010111000000100011100101";
wait for Clk_period;
Addr <= "0000111100000";
Trees_din <= "00000000000000110000100011100101";
wait for Clk_period;
Addr <= "0000111100001";
Trees_din <= "00000011000000000010111100000100";
wait for Clk_period;
Addr <= "0000111100010";
Trees_din <= "00000000001010110000100011100101";
wait for Clk_period;
Addr <= "0000111100011";
Trees_din <= "00000000001001010000100011100101";
wait for Clk_period;
Addr <= "0000111100100";
Trees_din <= "00000110000000000101000000001000";
wait for Clk_period;
Addr <= "0000111100101";
Trees_din <= "00000010000000000010111100000100";
wait for Clk_period;
Addr <= "0000111100110";
Trees_din <= "00000000010011110000100011100101";
wait for Clk_period;
Addr <= "0000111100111";
Trees_din <= "00000000000110100000100011100101";
wait for Clk_period;
Addr <= "0000111101000";
Trees_din <= "00000101000000000101100100000100";
wait for Clk_period;
Addr <= "0000111101001";
Trees_din <= "00000000000111010000100011100101";
wait for Clk_period;
Addr <= "0000111101010";
Trees_din <= "00000000010011000000100011100101";
wait for Clk_period;
Addr <= "0000111101011";
Trees_din <= "00000111000000000000111100010000";
wait for Clk_period;
Addr <= "0000111101100";
Trees_din <= "00000101000000000100110100001000";
wait for Clk_period;
Addr <= "0000111101101";
Trees_din <= "00000001000000000001000000000100";
wait for Clk_period;
Addr <= "0000111101110";
Trees_din <= "00000000001001110000100011100101";
wait for Clk_period;
Addr <= "0000111101111";
Trees_din <= "00000000010111100000100011100101";
wait for Clk_period;
Addr <= "0000111110000";
Trees_din <= "00000000000000000010011000000100";
wait for Clk_period;
Addr <= "0000111110001";
Trees_din <= "00000000000000110000100011100101";
wait for Clk_period;
Addr <= "0000111110010";
Trees_din <= "00000000000111010000100011100101";
wait for Clk_period;
Addr <= "0000111110011";
Trees_din <= "00000101000000000001111000001000";
wait for Clk_period;
Addr <= "0000111110100";
Trees_din <= "00000111000000000101011000000100";
wait for Clk_period;
Addr <= "0000111110101";
Trees_din <= "00000000001011000000100011100101";
wait for Clk_period;
Addr <= "0000111110110";
Trees_din <= "00000000001100010000100011100101";
wait for Clk_period;
Addr <= "0000111110111";
Trees_din <= "00000010000000000001011000000100";
wait for Clk_period;
Addr <= "0000111111000";
Trees_din <= "00000000010010110000100011100101";
wait for Clk_period;
Addr <= "0000111111001";
Trees_din <= "00000000000010010000100011100101";
wait for Clk_period;
Addr <= "0000111111010";
Trees_din <= "00000110000000000100000001000000";
wait for Clk_period;
Addr <= "0000111111011";
Trees_din <= "00000110000000000010001100100000";
wait for Clk_period;
Addr <= "0000111111100";
Trees_din <= "00000000000000000001000000010000";
wait for Clk_period;
Addr <= "0000111111101";
Trees_din <= "00000100000000000110000000001000";
wait for Clk_period;
Addr <= "0000111111110";
Trees_din <= "00000011000000000100100100000100";
wait for Clk_period;
Addr <= "0000111111111";
Trees_din <= "00000000010000000000100011100101";
wait for Clk_period;
Addr <= "0001000000000";
Trees_din <= "00000000010101010000100011100101";
wait for Clk_period;
Addr <= "0001000000001";
Trees_din <= "00000110000000000101111100000100";
wait for Clk_period;
Addr <= "0001000000010";
Trees_din <= "00000000001110110000100011100101";
wait for Clk_period;
Addr <= "0001000000011";
Trees_din <= "00000000001100110000100011100101";
wait for Clk_period;
Addr <= "0001000000100";
Trees_din <= "00000000000000000101001100001000";
wait for Clk_period;
Addr <= "0001000000101";
Trees_din <= "00000111000000000101101000000100";
wait for Clk_period;
Addr <= "0001000000110";
Trees_din <= "00000000000101010000100011100101";
wait for Clk_period;
Addr <= "0001000000111";
Trees_din <= "00000000010101100000100011100101";
wait for Clk_period;
Addr <= "0001000001000";
Trees_din <= "00000101000000000000000100000100";
wait for Clk_period;
Addr <= "0001000001001";
Trees_din <= "00000000000010010000100011100101";
wait for Clk_period;
Addr <= "0001000001010";
Trees_din <= "00000000000110000000100011100101";
wait for Clk_period;
Addr <= "0001000001011";
Trees_din <= "00000100000000000010111000010000";
wait for Clk_period;
Addr <= "0001000001100";
Trees_din <= "00000101000000000100000100001000";
wait for Clk_period;
Addr <= "0001000001101";
Trees_din <= "00000110000000000011110000000100";
wait for Clk_period;
Addr <= "0001000001110";
Trees_din <= "00000000000011100000100011100101";
wait for Clk_period;
Addr <= "0001000001111";
Trees_din <= "00000000000010000000100011100101";
wait for Clk_period;
Addr <= "0001000010000";
Trees_din <= "00000010000000000010110000000100";
wait for Clk_period;
Addr <= "0001000010001";
Trees_din <= "00000000000010000000100011100101";
wait for Clk_period;
Addr <= "0001000010010";
Trees_din <= "00000000001111000000100011100101";
wait for Clk_period;
Addr <= "0001000010011";
Trees_din <= "00000111000000000010000100001000";
wait for Clk_period;
Addr <= "0001000010100";
Trees_din <= "00000000000000000100011100000100";
wait for Clk_period;
Addr <= "0001000010101";
Trees_din <= "00000000000000110000100011100101";
wait for Clk_period;
Addr <= "0001000010110";
Trees_din <= "00000000000101100000100011100101";
wait for Clk_period;
Addr <= "0001000010111";
Trees_din <= "00000100000000000011100100000100";
wait for Clk_period;
Addr <= "0001000011000";
Trees_din <= "00000000000100010000100011100101";
wait for Clk_period;
Addr <= "0001000011001";
Trees_din <= "00000000000111000000100011100101";
wait for Clk_period;
Addr <= "0001000011010";
Trees_din <= "00000101000000000011100000100000";
wait for Clk_period;
Addr <= "0001000011011";
Trees_din <= "00000011000000000010000000010000";
wait for Clk_period;
Addr <= "0001000011100";
Trees_din <= "00000001000000000010111000001000";
wait for Clk_period;
Addr <= "0001000011101";
Trees_din <= "00000100000000000101010100000100";
wait for Clk_period;
Addr <= "0001000011110";
Trees_din <= "00000000001111100000100011100101";
wait for Clk_period;
Addr <= "0001000011111";
Trees_din <= "00000000000000100000100011100101";
wait for Clk_period;
Addr <= "0001000100000";
Trees_din <= "00000100000000000010000000000100";
wait for Clk_period;
Addr <= "0001000100001";
Trees_din <= "00000000001011010000100011100101";
wait for Clk_period;
Addr <= "0001000100010";
Trees_din <= "00000000001101010000100011100101";
wait for Clk_period;
Addr <= "0001000100011";
Trees_din <= "00000000000000000101111000001000";
wait for Clk_period;
Addr <= "0001000100100";
Trees_din <= "00000111000000000010001100000100";
wait for Clk_period;
Addr <= "0001000100101";
Trees_din <= "00000000001001000000100011100101";
wait for Clk_period;
Addr <= "0001000100110";
Trees_din <= "00000000001000000000100011100101";
wait for Clk_period;
Addr <= "0001000100111";
Trees_din <= "00000001000000000011001100000100";
wait for Clk_period;
Addr <= "0001000101000";
Trees_din <= "00000000000111100000100011100101";
wait for Clk_period;
Addr <= "0001000101001";
Trees_din <= "00000000000001110000100011100101";
wait for Clk_period;
Addr <= "0001000101010";
Trees_din <= "00000101000000000100100100010000";
wait for Clk_period;
Addr <= "0001000101011";
Trees_din <= "00000110000000000101010100001000";
wait for Clk_period;
Addr <= "0001000101100";
Trees_din <= "00000011000000000011010000000100";
wait for Clk_period;
Addr <= "0001000101101";
Trees_din <= "00000000000011110000100011100101";
wait for Clk_period;
Addr <= "0001000101110";
Trees_din <= "00000000001001100000100011100101";
wait for Clk_period;
Addr <= "0001000101111";
Trees_din <= "00000110000000000000101000000100";
wait for Clk_period;
Addr <= "0001000110000";
Trees_din <= "00000000000110110000100011100101";
wait for Clk_period;
Addr <= "0001000110001";
Trees_din <= "00000000001100100000100011100101";
wait for Clk_period;
Addr <= "0001000110010";
Trees_din <= "00000101000000000100101100001000";
wait for Clk_period;
Addr <= "0001000110011";
Trees_din <= "00000100000000000011000000000100";
wait for Clk_period;
Addr <= "0001000110100";
Trees_din <= "00000000001011100000100011100101";
wait for Clk_period;
Addr <= "0001000110101";
Trees_din <= "00000000000010010000100011100101";
wait for Clk_period;
Addr <= "0001000110110";
Trees_din <= "00000010000000000000110100000100";
wait for Clk_period;
Addr <= "0001000110111";
Trees_din <= "00000000001000010000100011100101";
wait for Clk_period;
Addr <= "0001000111000";
Trees_din <= "00000000010011110000100011100101";
wait for Clk_period;



----------tree 4-------------------

Addr <= "0001000111001";
Trees_din <= "00000000000000000010100010000000";
wait for Clk_period;
Addr <= "0001000111010";
Trees_din <= "00000101000000000011010101000000";
wait for Clk_period;
Addr <= "0001000111011";
Trees_din <= "00000110000000000010010000100000";
wait for Clk_period;
Addr <= "0001000111100";
Trees_din <= "00000001000000000101110100010000";
wait for Clk_period;
Addr <= "0001000111101";
Trees_din <= "00000111000000000001000100001000";
wait for Clk_period;
Addr <= "0001000111110";
Trees_din <= "00000000000000000010011100000100";
wait for Clk_period;
Addr <= "0001000111111";
Trees_din <= "00000000000001010000101011100001";
wait for Clk_period;
Addr <= "0001001000000";
Trees_din <= "00000000010100110000101011100001";
wait for Clk_period;
Addr <= "0001001000001";
Trees_din <= "00000000000000000001010100000100";
wait for Clk_period;
Addr <= "0001001000010";
Trees_din <= "00000000001011100000101011100001";
wait for Clk_period;
Addr <= "0001001000011";
Trees_din <= "00000000001000100000101011100001";
wait for Clk_period;
Addr <= "0001001000100";
Trees_din <= "00000001000000000100100000001000";
wait for Clk_period;
Addr <= "0001001000101";
Trees_din <= "00000101000000000000100100000100";
wait for Clk_period;
Addr <= "0001001000110";
Trees_din <= "00000000001111010000101011100001";
wait for Clk_period;
Addr <= "0001001000111";
Trees_din <= "00000000010001000000101011100001";
wait for Clk_period;
Addr <= "0001001001000";
Trees_din <= "00000000000000000011100100000100";
wait for Clk_period;
Addr <= "0001001001001";
Trees_din <= "00000000001001010000101011100001";
wait for Clk_period;
Addr <= "0001001001010";
Trees_din <= "00000000010101000000101011100001";
wait for Clk_period;
Addr <= "0001001001011";
Trees_din <= "00000010000000000101011100010000";
wait for Clk_period;
Addr <= "0001001001100";
Trees_din <= "00000110000000000011001100001000";
wait for Clk_period;
Addr <= "0001001001101";
Trees_din <= "00000010000000000010100000000100";
wait for Clk_period;
Addr <= "0001001001110";
Trees_din <= "00000000001101110000101011100001";
wait for Clk_period;
Addr <= "0001001001111";
Trees_din <= "00000000001000110000101011100001";
wait for Clk_period;
Addr <= "0001001010000";
Trees_din <= "00000100000000000100001100000100";
wait for Clk_period;
Addr <= "0001001010001";
Trees_din <= "00000000010110100000101011100001";
wait for Clk_period;
Addr <= "0001001010010";
Trees_din <= "00000000000100100000101011100001";
wait for Clk_period;
Addr <= "0001001010011";
Trees_din <= "00000110000000000000010100001000";
wait for Clk_period;
Addr <= "0001001010100";
Trees_din <= "00000100000000000000100100000100";
wait for Clk_period;
Addr <= "0001001010101";
Trees_din <= "00000000010111100000101011100001";
wait for Clk_period;
Addr <= "0001001010110";
Trees_din <= "00000000001110010000101011100001";
wait for Clk_period;
Addr <= "0001001010111";
Trees_din <= "00000111000000000100010000000100";
wait for Clk_period;
Addr <= "0001001011000";
Trees_din <= "00000000000101110000101011100001";
wait for Clk_period;
Addr <= "0001001011001";
Trees_din <= "00000000000110000000101011100001";
wait for Clk_period;
Addr <= "0001001011010";
Trees_din <= "00000011000000000100101000100000";
wait for Clk_period;
Addr <= "0001001011011";
Trees_din <= "00000100000000000011010100010000";
wait for Clk_period;
Addr <= "0001001011100";
Trees_din <= "00000111000000000000001000001000";
wait for Clk_period;
Addr <= "0001001011101";
Trees_din <= "00000011000000000001101000000100";
wait for Clk_period;
Addr <= "0001001011110";
Trees_din <= "00000000000010100000101011100001";
wait for Clk_period;
Addr <= "0001001011111";
Trees_din <= "00000000001001010000101011100001";
wait for Clk_period;
Addr <= "0001001100000";
Trees_din <= "00000100000000000010010100000100";
wait for Clk_period;
Addr <= "0001001100001";
Trees_din <= "00000000010100100000101011100001";
wait for Clk_period;
Addr <= "0001001100010";
Trees_din <= "00000000001000010000101011100001";
wait for Clk_period;
Addr <= "0001001100011";
Trees_din <= "00000000000000000001001000001000";
wait for Clk_period;
Addr <= "0001001100100";
Trees_din <= "00000100000000000101110100000100";
wait for Clk_period;
Addr <= "0001001100101";
Trees_din <= "00000000011001000000101011100001";
wait for Clk_period;
Addr <= "0001001100110";
Trees_din <= "00000000011001000000101011100001";
wait for Clk_period;
Addr <= "0001001100111";
Trees_din <= "00000001000000000110001000000100";
wait for Clk_period;
Addr <= "0001001101000";
Trees_din <= "00000000010000000000101011100001";
wait for Clk_period;
Addr <= "0001001101001";
Trees_din <= "00000000010110000000101011100001";
wait for Clk_period;
Addr <= "0001001101010";
Trees_din <= "00000100000000000001010100010000";
wait for Clk_period;
Addr <= "0001001101011";
Trees_din <= "00000100000000000010001100001000";
wait for Clk_period;
Addr <= "0001001101100";
Trees_din <= "00000101000000000101110100000100";
wait for Clk_period;
Addr <= "0001001101101";
Trees_din <= "00000000000101000000101011100001";
wait for Clk_period;
Addr <= "0001001101110";
Trees_din <= "00000000010110010000101011100001";
wait for Clk_period;
Addr <= "0001001101111";
Trees_din <= "00000101000000000011100100000100";
wait for Clk_period;
Addr <= "0001001110000";
Trees_din <= "00000000011000000000101011100001";
wait for Clk_period;
Addr <= "0001001110001";
Trees_din <= "00000000000100010000101011100001";
wait for Clk_period;
Addr <= "0001001110010";
Trees_din <= "00000011000000000011101000001000";
wait for Clk_period;
Addr <= "0001001110011";
Trees_din <= "00000111000000000001011000000100";
wait for Clk_period;
Addr <= "0001001110100";
Trees_din <= "00000000001100010000101011100001";
wait for Clk_period;
Addr <= "0001001110101";
Trees_din <= "00000000000111010000101011100001";
wait for Clk_period;
Addr <= "0001001110110";
Trees_din <= "00000110000000000101100100000100";
wait for Clk_period;
Addr <= "0001001110111";
Trees_din <= "00000000010000110000101011100001";
wait for Clk_period;
Addr <= "0001001111000";
Trees_din <= "00000000000111100000101011100001";
wait for Clk_period;
Addr <= "0001001111001";
Trees_din <= "00000100000000000100111001000000";
wait for Clk_period;
Addr <= "0001001111010";
Trees_din <= "00000011000000000110001000100000";
wait for Clk_period;
Addr <= "0001001111011";
Trees_din <= "00000011000000000010001000010000";
wait for Clk_period;
Addr <= "0001001111100";
Trees_din <= "00000011000000000001100100001000";
wait for Clk_period;
Addr <= "0001001111101";
Trees_din <= "00000110000000000011101100000100";
wait for Clk_period;
Addr <= "0001001111110";
Trees_din <= "00000000010110000000101011100001";
wait for Clk_period;
Addr <= "0001001111111";
Trees_din <= "00000000001001110000101011100001";
wait for Clk_period;
Addr <= "0001010000000";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0001010000001";
Trees_din <= "00000000010010010000101011100001";
wait for Clk_period;
Addr <= "0001010000010";
Trees_din <= "00000000000000110000101011100001";
wait for Clk_period;
Addr <= "0001010000011";
Trees_din <= "00000001000000000101010000001000";
wait for Clk_period;
Addr <= "0001010000100";
Trees_din <= "00000111000000000100010100000100";
wait for Clk_period;
Addr <= "0001010000101";
Trees_din <= "00000000010011010000101011100001";
wait for Clk_period;
Addr <= "0001010000110";
Trees_din <= "00000000001011000000101011100001";
wait for Clk_period;
Addr <= "0001010000111";
Trees_din <= "00000101000000000000001000000100";
wait for Clk_period;
Addr <= "0001010001000";
Trees_din <= "00000000010010110000101011100001";
wait for Clk_period;
Addr <= "0001010001001";
Trees_din <= "00000000000000100000101011100001";
wait for Clk_period;
Addr <= "0001010001010";
Trees_din <= "00000110000000000100100000010000";
wait for Clk_period;
Addr <= "0001010001011";
Trees_din <= "00000101000000000010101100001000";
wait for Clk_period;
Addr <= "0001010001100";
Trees_din <= "00000100000000000001110000000100";
wait for Clk_period;
Addr <= "0001010001101";
Trees_din <= "00000000001110110000101011100001";
wait for Clk_period;
Addr <= "0001010001110";
Trees_din <= "00000000010000010000101011100001";
wait for Clk_period;
Addr <= "0001010001111";
Trees_din <= "00000001000000000100101000000100";
wait for Clk_period;
Addr <= "0001010010000";
Trees_din <= "00000000010001100000101011100001";
wait for Clk_period;
Addr <= "0001010010001";
Trees_din <= "00000000001110100000101011100001";
wait for Clk_period;
Addr <= "0001010010010";
Trees_din <= "00000011000000000000010000001000";
wait for Clk_period;
Addr <= "0001010010011";
Trees_din <= "00000000000000000010100000000100";
wait for Clk_period;
Addr <= "0001010010100";
Trees_din <= "00000000000011100000101011100001";
wait for Clk_period;
Addr <= "0001010010101";
Trees_din <= "00000000011000100000101011100001";
wait for Clk_period;
Addr <= "0001010010110";
Trees_din <= "00000100000000000000111000000100";
wait for Clk_period;
Addr <= "0001010010111";
Trees_din <= "00000000000011000000101011100001";
wait for Clk_period;
Addr <= "0001010011000";
Trees_din <= "00000000010010010000101011100001";
wait for Clk_period;
Addr <= "0001010011001";
Trees_din <= "00000101000000000010010000100000";
wait for Clk_period;
Addr <= "0001010011010";
Trees_din <= "00000000000000000101000000010000";
wait for Clk_period;
Addr <= "0001010011011";
Trees_din <= "00000010000000000101001100001000";
wait for Clk_period;
Addr <= "0001010011100";
Trees_din <= "00000010000000000100010100000100";
wait for Clk_period;
Addr <= "0001010011101";
Trees_din <= "00000000001001000000101011100001";
wait for Clk_period;
Addr <= "0001010011110";
Trees_din <= "00000000001100000000101011100001";
wait for Clk_period;
Addr <= "0001010011111";
Trees_din <= "00000000000000000000010000000100";
wait for Clk_period;
Addr <= "0001010100000";
Trees_din <= "00000000001110000000101011100001";
wait for Clk_period;
Addr <= "0001010100001";
Trees_din <= "00000000000000010000101011100001";
wait for Clk_period;
Addr <= "0001010100010";
Trees_din <= "00000000000000000011111000001000";
wait for Clk_period;
Addr <= "0001010100011";
Trees_din <= "00000000000000000010000100000100";
wait for Clk_period;
Addr <= "0001010100100";
Trees_din <= "00000000010000010000101011100001";
wait for Clk_period;
Addr <= "0001010100101";
Trees_din <= "00000000000100000000101011100001";
wait for Clk_period;
Addr <= "0001010100110";
Trees_din <= "00000100000000000101110100000100";
wait for Clk_period;
Addr <= "0001010100111";
Trees_din <= "00000000000011110000101011100001";
wait for Clk_period;
Addr <= "0001010101000";
Trees_din <= "00000000001001110000101011100001";
wait for Clk_period;
Addr <= "0001010101001";
Trees_din <= "00000110000000000010000100010000";
wait for Clk_period;
Addr <= "0001010101010";
Trees_din <= "00000011000000000000010000001000";
wait for Clk_period;
Addr <= "0001010101011";
Trees_din <= "00000010000000000101100000000100";
wait for Clk_period;
Addr <= "0001010101100";
Trees_din <= "00000000000111100000101011100001";
wait for Clk_period;
Addr <= "0001010101101";
Trees_din <= "00000000001110100000101011100001";
wait for Clk_period;
Addr <= "0001010101110";
Trees_din <= "00000000000000000010010000000100";
wait for Clk_period;
Addr <= "0001010101111";
Trees_din <= "00000000000110010000101011100001";
wait for Clk_period;
Addr <= "0001010110000";
Trees_din <= "00000000010010010000101011100001";
wait for Clk_period;
Addr <= "0001010110001";
Trees_din <= "00000111000000000011111100001000";
wait for Clk_period;
Addr <= "0001010110010";
Trees_din <= "00000010000000000001001100000100";
wait for Clk_period;
Addr <= "0001010110011";
Trees_din <= "00000000001111110000101011100001";
wait for Clk_period;
Addr <= "0001010110100";
Trees_din <= "00000000000101000000101011100001";
wait for Clk_period;
Addr <= "0001010110101";
Trees_din <= "00000001000000000011011100000100";
wait for Clk_period;
Addr <= "0001010110110";
Trees_din <= "00000000000000100000101011100001";
wait for Clk_period;
Addr <= "0001010110111";
Trees_din <= "00000000010001010000101011100001";
wait for Clk_period;



----------tree 5-------------------

Addr <= "0001010111000";
Trees_din <= "00000100000000000000001110000000";
wait for Clk_period;
Addr <= "0001010111001";
Trees_din <= "00000100000000000011100101000000";
wait for Clk_period;
Addr <= "0001010111010";
Trees_din <= "00000110000000000110000000100000";
wait for Clk_period;
Addr <= "0001010111011";
Trees_din <= "00000111000000000000101000010000";
wait for Clk_period;
Addr <= "0001010111100";
Trees_din <= "00000001000000000100111100001000";
wait for Clk_period;
Addr <= "0001010111101";
Trees_din <= "00000100000000000100001100000100";
wait for Clk_period;
Addr <= "0001010111110";
Trees_din <= "00000000001000000000110011011101";
wait for Clk_period;
Addr <= "0001010111111";
Trees_din <= "00000000001001010000110011011101";
wait for Clk_period;
Addr <= "0001011000000";
Trees_din <= "00000000000000000011111000000100";
wait for Clk_period;
Addr <= "0001011000001";
Trees_din <= "00000000001100110000110011011101";
wait for Clk_period;
Addr <= "0001011000010";
Trees_din <= "00000000000110010000110011011101";
wait for Clk_period;
Addr <= "0001011000011";
Trees_din <= "00000001000000000001111100001000";
wait for Clk_period;
Addr <= "0001011000100";
Trees_din <= "00000101000000000110010000000100";
wait for Clk_period;
Addr <= "0001011000101";
Trees_din <= "00000000000010110000110011011101";
wait for Clk_period;
Addr <= "0001011000110";
Trees_din <= "00000000000101000000110011011101";
wait for Clk_period;
Addr <= "0001011000111";
Trees_din <= "00000101000000000000111100000100";
wait for Clk_period;
Addr <= "0001011001000";
Trees_din <= "00000000001001110000110011011101";
wait for Clk_period;
Addr <= "0001011001001";
Trees_din <= "00000000000001000000110011011101";
wait for Clk_period;
Addr <= "0001011001010";
Trees_din <= "00000000000000000101000100010000";
wait for Clk_period;
Addr <= "0001011001011";
Trees_din <= "00000111000000000101100000001000";
wait for Clk_period;
Addr <= "0001011001100";
Trees_din <= "00000001000000000010101000000100";
wait for Clk_period;
Addr <= "0001011001101";
Trees_din <= "00000000010111000000110011011101";
wait for Clk_period;
Addr <= "0001011001110";
Trees_din <= "00000000000011010000110011011101";
wait for Clk_period;
Addr <= "0001011001111";
Trees_din <= "00000101000000000000110100000100";
wait for Clk_period;
Addr <= "0001011010000";
Trees_din <= "00000000001111110000110011011101";
wait for Clk_period;
Addr <= "0001011010001";
Trees_din <= "00000000001110110000110011011101";
wait for Clk_period;
Addr <= "0001011010010";
Trees_din <= "00000101000000000001001100001000";
wait for Clk_period;
Addr <= "0001011010011";
Trees_din <= "00000110000000000000101000000100";
wait for Clk_period;
Addr <= "0001011010100";
Trees_din <= "00000000010001010000110011011101";
wait for Clk_period;
Addr <= "0001011010101";
Trees_din <= "00000000010100110000110011011101";
wait for Clk_period;
Addr <= "0001011010110";
Trees_din <= "00000000000000000001010000000100";
wait for Clk_period;
Addr <= "0001011010111";
Trees_din <= "00000000011000100000110011011101";
wait for Clk_period;
Addr <= "0001011011000";
Trees_din <= "00000000001111000000110011011101";
wait for Clk_period;
Addr <= "0001011011001";
Trees_din <= "00000111000000000010100100100000";
wait for Clk_period;
Addr <= "0001011011010";
Trees_din <= "00000111000000000000100100010000";
wait for Clk_period;
Addr <= "0001011011011";
Trees_din <= "00000110000000000010101000001000";
wait for Clk_period;
Addr <= "0001011011100";
Trees_din <= "00000011000000000010011000000100";
wait for Clk_period;
Addr <= "0001011011101";
Trees_din <= "00000000001000110000110011011101";
wait for Clk_period;
Addr <= "0001011011110";
Trees_din <= "00000000000010010000110011011101";
wait for Clk_period;
Addr <= "0001011011111";
Trees_din <= "00000100000000000001111000000100";
wait for Clk_period;
Addr <= "0001011100000";
Trees_din <= "00000000010000010000110011011101";
wait for Clk_period;
Addr <= "0001011100001";
Trees_din <= "00000000000101010000110011011101";
wait for Clk_period;
Addr <= "0001011100010";
Trees_din <= "00000010000000000010010100001000";
wait for Clk_period;
Addr <= "0001011100011";
Trees_din <= "00000000000000000011111100000100";
wait for Clk_period;
Addr <= "0001011100100";
Trees_din <= "00000000000100110000110011011101";
wait for Clk_period;
Addr <= "0001011100101";
Trees_din <= "00000000001011100000110011011101";
wait for Clk_period;
Addr <= "0001011100110";
Trees_din <= "00000011000000000000101100000100";
wait for Clk_period;
Addr <= "0001011100111";
Trees_din <= "00000000010110000000110011011101";
wait for Clk_period;
Addr <= "0001011101000";
Trees_din <= "00000000000110000000110011011101";
wait for Clk_period;
Addr <= "0001011101001";
Trees_din <= "00000011000000000001011000010000";
wait for Clk_period;
Addr <= "0001011101010";
Trees_din <= "00000101000000000100110100001000";
wait for Clk_period;
Addr <= "0001011101011";
Trees_din <= "00000101000000000110001100000100";
wait for Clk_period;
Addr <= "0001011101100";
Trees_din <= "00000000000000110000110011011101";
wait for Clk_period;
Addr <= "0001011101101";
Trees_din <= "00000000000011000000110011011101";
wait for Clk_period;
Addr <= "0001011101110";
Trees_din <= "00000001000000000011011100000100";
wait for Clk_period;
Addr <= "0001011101111";
Trees_din <= "00000000000011000000110011011101";
wait for Clk_period;
Addr <= "0001011110000";
Trees_din <= "00000000001101010000110011011101";
wait for Clk_period;
Addr <= "0001011110001";
Trees_din <= "00000100000000000101001000001000";
wait for Clk_period;
Addr <= "0001011110010";
Trees_din <= "00000000000000000100010000000100";
wait for Clk_period;
Addr <= "0001011110011";
Trees_din <= "00000000010010100000110011011101";
wait for Clk_period;
Addr <= "0001011110100";
Trees_din <= "00000000010000010000110011011101";
wait for Clk_period;
Addr <= "0001011110101";
Trees_din <= "00000111000000000000101100000100";
wait for Clk_period;
Addr <= "0001011110110";
Trees_din <= "00000000001110110000110011011101";
wait for Clk_period;
Addr <= "0001011110111";
Trees_din <= "00000000010101010000110011011101";
wait for Clk_period;
Addr <= "0001011111000";
Trees_din <= "00000010000000000000110101000000";
wait for Clk_period;
Addr <= "0001011111001";
Trees_din <= "00000010000000000001000000100000";
wait for Clk_period;
Addr <= "0001011111010";
Trees_din <= "00000110000000000001011100010000";
wait for Clk_period;
Addr <= "0001011111011";
Trees_din <= "00000110000000000100011000001000";
wait for Clk_period;
Addr <= "0001011111100";
Trees_din <= "00000110000000000110001000000100";
wait for Clk_period;
Addr <= "0001011111101";
Trees_din <= "00000000000101010000110011011101";
wait for Clk_period;
Addr <= "0001011111110";
Trees_din <= "00000000000101010000110011011101";
wait for Clk_period;
Addr <= "0001011111111";
Trees_din <= "00000101000000000000001000000100";
wait for Clk_period;
Addr <= "0001100000000";
Trees_din <= "00000000000010010000110011011101";
wait for Clk_period;
Addr <= "0001100000001";
Trees_din <= "00000000001101100000110011011101";
wait for Clk_period;
Addr <= "0001100000010";
Trees_din <= "00000111000000000010000000001000";
wait for Clk_period;
Addr <= "0001100000011";
Trees_din <= "00000110000000000001101100000100";
wait for Clk_period;
Addr <= "0001100000100";
Trees_din <= "00000000000110100000110011011101";
wait for Clk_period;
Addr <= "0001100000101";
Trees_din <= "00000000010001010000110011011101";
wait for Clk_period;
Addr <= "0001100000110";
Trees_din <= "00000010000000000000111100000100";
wait for Clk_period;
Addr <= "0001100000111";
Trees_din <= "00000000010110000000110011011101";
wait for Clk_period;
Addr <= "0001100001000";
Trees_din <= "00000000010101110000110011011101";
wait for Clk_period;
Addr <= "0001100001001";
Trees_din <= "00000110000000000101000100010000";
wait for Clk_period;
Addr <= "0001100001010";
Trees_din <= "00000010000000000010000000001000";
wait for Clk_period;
Addr <= "0001100001011";
Trees_din <= "00000011000000000011110100000100";
wait for Clk_period;
Addr <= "0001100001100";
Trees_din <= "00000000000011100000110011011101";
wait for Clk_period;
Addr <= "0001100001101";
Trees_din <= "00000000001111010000110011011101";
wait for Clk_period;
Addr <= "0001100001110";
Trees_din <= "00000010000000000010000100000100";
wait for Clk_period;
Addr <= "0001100001111";
Trees_din <= "00000000000011110000110011011101";
wait for Clk_period;
Addr <= "0001100010000";
Trees_din <= "00000000001000100000110011011101";
wait for Clk_period;
Addr <= "0001100010001";
Trees_din <= "00000000000000000000011100001000";
wait for Clk_period;
Addr <= "0001100010010";
Trees_din <= "00000010000000000000000100000100";
wait for Clk_period;
Addr <= "0001100010011";
Trees_din <= "00000000010001010000110011011101";
wait for Clk_period;
Addr <= "0001100010100";
Trees_din <= "00000000001001010000110011011101";
wait for Clk_period;
Addr <= "0001100010101";
Trees_din <= "00000101000000000001100000000100";
wait for Clk_period;
Addr <= "0001100010110";
Trees_din <= "00000000010011100000110011011101";
wait for Clk_period;
Addr <= "0001100010111";
Trees_din <= "00000000001100110000110011011101";
wait for Clk_period;
Addr <= "0001100011000";
Trees_din <= "00000011000000000001011100100000";
wait for Clk_period;
Addr <= "0001100011001";
Trees_din <= "00000110000000000001010100010000";
wait for Clk_period;
Addr <= "0001100011010";
Trees_din <= "00000110000000000000101100001000";
wait for Clk_period;
Addr <= "0001100011011";
Trees_din <= "00000111000000000001001000000100";
wait for Clk_period;
Addr <= "0001100011100";
Trees_din <= "00000000010111000000110011011101";
wait for Clk_period;
Addr <= "0001100011101";
Trees_din <= "00000000001100010000110011011101";
wait for Clk_period;
Addr <= "0001100011110";
Trees_din <= "00000001000000000000011100000100";
wait for Clk_period;
Addr <= "0001100011111";
Trees_din <= "00000000011000000000110011011101";
wait for Clk_period;
Addr <= "0001100100000";
Trees_din <= "00000000010111110000110011011101";
wait for Clk_period;
Addr <= "0001100100001";
Trees_din <= "00000001000000000010101100001000";
wait for Clk_period;
Addr <= "0001100100010";
Trees_din <= "00000111000000000011100000000100";
wait for Clk_period;
Addr <= "0001100100011";
Trees_din <= "00000000010000010000110011011101";
wait for Clk_period;
Addr <= "0001100100100";
Trees_din <= "00000000000001110000110011011101";
wait for Clk_period;
Addr <= "0001100100101";
Trees_din <= "00000011000000000101001100000100";
wait for Clk_period;
Addr <= "0001100100110";
Trees_din <= "00000000010010110000110011011101";
wait for Clk_period;
Addr <= "0001100100111";
Trees_din <= "00000000000110100000110011011101";
wait for Clk_period;
Addr <= "0001100101000";
Trees_din <= "00000100000000000000001000010000";
wait for Clk_period;
Addr <= "0001100101001";
Trees_din <= "00000001000000000010010000001000";
wait for Clk_period;
Addr <= "0001100101010";
Trees_din <= "00000010000000000001110100000100";
wait for Clk_period;
Addr <= "0001100101011";
Trees_din <= "00000000010101010000110011011101";
wait for Clk_period;
Addr <= "0001100101100";
Trees_din <= "00000000010110000000110011011101";
wait for Clk_period;
Addr <= "0001100101101";
Trees_din <= "00000001000000000010111100000100";
wait for Clk_period;
Addr <= "0001100101110";
Trees_din <= "00000000010000010000110011011101";
wait for Clk_period;
Addr <= "0001100101111";
Trees_din <= "00000000000110100000110011011101";
wait for Clk_period;
Addr <= "0001100110000";
Trees_din <= "00000001000000000011011000001000";
wait for Clk_period;
Addr <= "0001100110001";
Trees_din <= "00000101000000000000111000000100";
wait for Clk_period;
Addr <= "0001100110010";
Trees_din <= "00000000000111000000110011011101";
wait for Clk_period;
Addr <= "0001100110011";
Trees_din <= "00000000000111110000110011011101";
wait for Clk_period;
Addr <= "0001100110100";
Trees_din <= "00000111000000000101111100000100";
wait for Clk_period;
Addr <= "0001100110101";
Trees_din <= "00000000011000010000110011011101";
wait for Clk_period;
Addr <= "0001100110110";
Trees_din <= "00000000001011110000110011011101";
wait for Clk_period;



----------tree 6-------------------

Addr <= "0001100110111";
Trees_din <= "00000010000000000100000110000000";
wait for Clk_period;
Addr <= "0001100111000";
Trees_din <= "00000111000000000101000101000000";
wait for Clk_period;
Addr <= "0001100111001";
Trees_din <= "00000001000000000010100100100000";
wait for Clk_period;
Addr <= "0001100111010";
Trees_din <= "00000111000000000101001000010000";
wait for Clk_period;
Addr <= "0001100111011";
Trees_din <= "00000001000000000101001000001000";
wait for Clk_period;
Addr <= "0001100111100";
Trees_din <= "00000000000000000010010100000100";
wait for Clk_period;
Addr <= "0001100111101";
Trees_din <= "00000000010001000000111011011001";
wait for Clk_period;
Addr <= "0001100111110";
Trees_din <= "00000000001101100000111011011001";
wait for Clk_period;
Addr <= "0001100111111";
Trees_din <= "00000111000000000001000000000100";
wait for Clk_period;
Addr <= "0001101000000";
Trees_din <= "00000000000100010000111011011001";
wait for Clk_period;
Addr <= "0001101000001";
Trees_din <= "00000000001111100000111011011001";
wait for Clk_period;
Addr <= "0001101000010";
Trees_din <= "00000110000000000010000000001000";
wait for Clk_period;
Addr <= "0001101000011";
Trees_din <= "00000101000000000011000000000100";
wait for Clk_period;
Addr <= "0001101000100";
Trees_din <= "00000000010110110000111011011001";
wait for Clk_period;
Addr <= "0001101000101";
Trees_din <= "00000000001110110000111011011001";
wait for Clk_period;
Addr <= "0001101000110";
Trees_din <= "00000100000000000010011000000100";
wait for Clk_period;
Addr <= "0001101000111";
Trees_din <= "00000000000100110000111011011001";
wait for Clk_period;
Addr <= "0001101001000";
Trees_din <= "00000000000111100000111011011001";
wait for Clk_period;
Addr <= "0001101001001";
Trees_din <= "00000100000000000101010100010000";
wait for Clk_period;
Addr <= "0001101001010";
Trees_din <= "00000100000000000000011100001000";
wait for Clk_period;
Addr <= "0001101001011";
Trees_din <= "00000000000000000001110000000100";
wait for Clk_period;
Addr <= "0001101001100";
Trees_din <= "00000000000111110000111011011001";
wait for Clk_period;
Addr <= "0001101001101";
Trees_din <= "00000000010010110000111011011001";
wait for Clk_period;
Addr <= "0001101001110";
Trees_din <= "00000110000000000010100000000100";
wait for Clk_period;
Addr <= "0001101001111";
Trees_din <= "00000000010111100000111011011001";
wait for Clk_period;
Addr <= "0001101010000";
Trees_din <= "00000000010100100000111011011001";
wait for Clk_period;
Addr <= "0001101010001";
Trees_din <= "00000011000000000010101100001000";
wait for Clk_period;
Addr <= "0001101010010";
Trees_din <= "00000011000000000101010000000100";
wait for Clk_period;
Addr <= "0001101010011";
Trees_din <= "00000000001110100000111011011001";
wait for Clk_period;
Addr <= "0001101010100";
Trees_din <= "00000000000101110000111011011001";
wait for Clk_period;
Addr <= "0001101010101";
Trees_din <= "00000001000000000001110000000100";
wait for Clk_period;
Addr <= "0001101010110";
Trees_din <= "00000000000011000000111011011001";
wait for Clk_period;
Addr <= "0001101010111";
Trees_din <= "00000000001001110000111011011001";
wait for Clk_period;
Addr <= "0001101011000";
Trees_din <= "00000000000000000101100000100000";
wait for Clk_period;
Addr <= "0001101011001";
Trees_din <= "00000001000000000000110000010000";
wait for Clk_period;
Addr <= "0001101011010";
Trees_din <= "00000011000000000100011100001000";
wait for Clk_period;
Addr <= "0001101011011";
Trees_din <= "00000101000000000100100000000100";
wait for Clk_period;
Addr <= "0001101011100";
Trees_din <= "00000000001000010000111011011001";
wait for Clk_period;
Addr <= "0001101011101";
Trees_din <= "00000000010000010000111011011001";
wait for Clk_period;
Addr <= "0001101011110";
Trees_din <= "00000011000000000101011000000100";
wait for Clk_period;
Addr <= "0001101011111";
Trees_din <= "00000000010111010000111011011001";
wait for Clk_period;
Addr <= "0001101100000";
Trees_din <= "00000000001011110000111011011001";
wait for Clk_period;
Addr <= "0001101100001";
Trees_din <= "00000011000000000001101100001000";
wait for Clk_period;
Addr <= "0001101100010";
Trees_din <= "00000111000000000001001000000100";
wait for Clk_period;
Addr <= "0001101100011";
Trees_din <= "00000000001000110000111011011001";
wait for Clk_period;
Addr <= "0001101100100";
Trees_din <= "00000000010101010000111011011001";
wait for Clk_period;
Addr <= "0001101100101";
Trees_din <= "00000010000000000001101100000100";
wait for Clk_period;
Addr <= "0001101100110";
Trees_din <= "00000000001111110000111011011001";
wait for Clk_period;
Addr <= "0001101100111";
Trees_din <= "00000000010011010000111011011001";
wait for Clk_period;
Addr <= "0001101101000";
Trees_din <= "00000110000000000101111100010000";
wait for Clk_period;
Addr <= "0001101101001";
Trees_din <= "00000100000000000001100100001000";
wait for Clk_period;
Addr <= "0001101101010";
Trees_din <= "00000001000000000010010100000100";
wait for Clk_period;
Addr <= "0001101101011";
Trees_din <= "00000000001001000000111011011001";
wait for Clk_period;
Addr <= "0001101101100";
Trees_din <= "00000000010101010000111011011001";
wait for Clk_period;
Addr <= "0001101101101";
Trees_din <= "00000001000000000000111000000100";
wait for Clk_period;
Addr <= "0001101101110";
Trees_din <= "00000000010110100000111011011001";
wait for Clk_period;
Addr <= "0001101101111";
Trees_din <= "00000000001100110000111011011001";
wait for Clk_period;
Addr <= "0001101110000";
Trees_din <= "00000001000000000001001100001000";
wait for Clk_period;
Addr <= "0001101110001";
Trees_din <= "00000001000000000000000100000100";
wait for Clk_period;
Addr <= "0001101110010";
Trees_din <= "00000000010010000000111011011001";
wait for Clk_period;
Addr <= "0001101110011";
Trees_din <= "00000000000001000000111011011001";
wait for Clk_period;
Addr <= "0001101110100";
Trees_din <= "00000100000000000101100000000100";
wait for Clk_period;
Addr <= "0001101110101";
Trees_din <= "00000000000010110000111011011001";
wait for Clk_period;
Addr <= "0001101110110";
Trees_din <= "00000000001111110000111011011001";
wait for Clk_period;
Addr <= "0001101110111";
Trees_din <= "00000010000000000011010001000000";
wait for Clk_period;
Addr <= "0001101111000";
Trees_din <= "00000000000000000100100100100000";
wait for Clk_period;
Addr <= "0001101111001";
Trees_din <= "00000100000000000010100000010000";
wait for Clk_period;
Addr <= "0001101111010";
Trees_din <= "00000010000000000101010100001000";
wait for Clk_period;
Addr <= "0001101111011";
Trees_din <= "00000010000000000011001100000100";
wait for Clk_period;
Addr <= "0001101111100";
Trees_din <= "00000000000000100000111011011001";
wait for Clk_period;
Addr <= "0001101111101";
Trees_din <= "00000000010100000000111011011001";
wait for Clk_period;
Addr <= "0001101111110";
Trees_din <= "00000110000000000000111000000100";
wait for Clk_period;
Addr <= "0001101111111";
Trees_din <= "00000000001000000000111011011001";
wait for Clk_period;
Addr <= "0001110000000";
Trees_din <= "00000000010001010000111011011001";
wait for Clk_period;
Addr <= "0001110000001";
Trees_din <= "00000111000000000000101000001000";
wait for Clk_period;
Addr <= "0001110000010";
Trees_din <= "00000010000000000011101000000100";
wait for Clk_period;
Addr <= "0001110000011";
Trees_din <= "00000000010001100000111011011001";
wait for Clk_period;
Addr <= "0001110000100";
Trees_din <= "00000000000111110000111011011001";
wait for Clk_period;
Addr <= "0001110000101";
Trees_din <= "00000001000000000101011000000100";
wait for Clk_period;
Addr <= "0001110000110";
Trees_din <= "00000000010001010000111011011001";
wait for Clk_period;
Addr <= "0001110000111";
Trees_din <= "00000000001000110000111011011001";
wait for Clk_period;
Addr <= "0001110001000";
Trees_din <= "00000000000000000010001100010000";
wait for Clk_period;
Addr <= "0001110001001";
Trees_din <= "00000100000000000011011100001000";
wait for Clk_period;
Addr <= "0001110001010";
Trees_din <= "00000110000000000101001000000100";
wait for Clk_period;
Addr <= "0001110001011";
Trees_din <= "00000000001111000000111011011001";
wait for Clk_period;
Addr <= "0001110001100";
Trees_din <= "00000000010001100000111011011001";
wait for Clk_period;
Addr <= "0001110001101";
Trees_din <= "00000111000000000101101100000100";
wait for Clk_period;
Addr <= "0001110001110";
Trees_din <= "00000000010110000000111011011001";
wait for Clk_period;
Addr <= "0001110001111";
Trees_din <= "00000000000110110000111011011001";
wait for Clk_period;
Addr <= "0001110010000";
Trees_din <= "00000101000000000100110000001000";
wait for Clk_period;
Addr <= "0001110010001";
Trees_din <= "00000000000000000100001100000100";
wait for Clk_period;
Addr <= "0001110010010";
Trees_din <= "00000000010001110000111011011001";
wait for Clk_period;
Addr <= "0001110010011";
Trees_din <= "00000000010111100000111011011001";
wait for Clk_period;
Addr <= "0001110010100";
Trees_din <= "00000011000000000000000100000100";
wait for Clk_period;
Addr <= "0001110010101";
Trees_din <= "00000000001010110000111011011001";
wait for Clk_period;
Addr <= "0001110010110";
Trees_din <= "00000000001000010000111011011001";
wait for Clk_period;
Addr <= "0001110010111";
Trees_din <= "00000110000000000011000000100000";
wait for Clk_period;
Addr <= "0001110011000";
Trees_din <= "00000111000000000110000100010000";
wait for Clk_period;
Addr <= "0001110011001";
Trees_din <= "00000111000000000100100100001000";
wait for Clk_period;
Addr <= "0001110011010";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "0001110011011";
Trees_din <= "00000000001001000000111011011001";
wait for Clk_period;
Addr <= "0001110011100";
Trees_din <= "00000000001110010000111011011001";
wait for Clk_period;
Addr <= "0001110011101";
Trees_din <= "00000011000000000010101100000100";
wait for Clk_period;
Addr <= "0001110011110";
Trees_din <= "00000000000101100000111011011001";
wait for Clk_period;
Addr <= "0001110011111";
Trees_din <= "00000000000000010000111011011001";
wait for Clk_period;
Addr <= "0001110100000";
Trees_din <= "00000010000000000100100100001000";
wait for Clk_period;
Addr <= "0001110100001";
Trees_din <= "00000110000000000010010000000100";
wait for Clk_period;
Addr <= "0001110100010";
Trees_din <= "00000000010001110000111011011001";
wait for Clk_period;
Addr <= "0001110100011";
Trees_din <= "00000000001111000000111011011001";
wait for Clk_period;
Addr <= "0001110100100";
Trees_din <= "00000101000000000011101000000100";
wait for Clk_period;
Addr <= "0001110100101";
Trees_din <= "00000000010011110000111011011001";
wait for Clk_period;
Addr <= "0001110100110";
Trees_din <= "00000000010001010000111011011001";
wait for Clk_period;
Addr <= "0001110100111";
Trees_din <= "00000111000000000010111100010000";
wait for Clk_period;
Addr <= "0001110101000";
Trees_din <= "00000011000000000011100000001000";
wait for Clk_period;
Addr <= "0001110101001";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "0001110101010";
Trees_din <= "00000000000000000000111011011001";
wait for Clk_period;
Addr <= "0001110101011";
Trees_din <= "00000000001001110000111011011001";
wait for Clk_period;
Addr <= "0001110101100";
Trees_din <= "00000001000000000001110000000100";
wait for Clk_period;
Addr <= "0001110101101";
Trees_din <= "00000000010101010000111011011001";
wait for Clk_period;
Addr <= "0001110101110";
Trees_din <= "00000000000000100000111011011001";
wait for Clk_period;
Addr <= "0001110101111";
Trees_din <= "00000111000000000100100000001000";
wait for Clk_period;
Addr <= "0001110110000";
Trees_din <= "00000110000000000100110100000100";
wait for Clk_period;
Addr <= "0001110110001";
Trees_din <= "00000000000001110000111011011001";
wait for Clk_period;
Addr <= "0001110110010";
Trees_din <= "00000000010001000000111011011001";
wait for Clk_period;
Addr <= "0001110110011";
Trees_din <= "00000100000000000000010100000100";
wait for Clk_period;
Addr <= "0001110110100";
Trees_din <= "00000000000110010000111011011001";
wait for Clk_period;
Addr <= "0001110110101";
Trees_din <= "00000000011000000000111011011001";
wait for Clk_period;



----------tree 7-------------------

Addr <= "0001110110110";
Trees_din <= "00000011000000000010110110000000";
wait for Clk_period;
Addr <= "0001110110111";
Trees_din <= "00000100000000000101101101000000";
wait for Clk_period;
Addr <= "0001110111000";
Trees_din <= "00000110000000000010001100100000";
wait for Clk_period;
Addr <= "0001110111001";
Trees_din <= "00000101000000000100011100010000";
wait for Clk_period;
Addr <= "0001110111010";
Trees_din <= "00000110000000000011010000001000";
wait for Clk_period;
Addr <= "0001110111011";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0001110111100";
Trees_din <= "00000000000100100001000011010101";
wait for Clk_period;
Addr <= "0001110111101";
Trees_din <= "00000000010100010001000011010101";
wait for Clk_period;
Addr <= "0001110111110";
Trees_din <= "00000111000000000000100100000100";
wait for Clk_period;
Addr <= "0001110111111";
Trees_din <= "00000000001001100001000011010101";
wait for Clk_period;
Addr <= "0001111000000";
Trees_din <= "00000000011001000001000011010101";
wait for Clk_period;
Addr <= "0001111000001";
Trees_din <= "00000001000000000000101000001000";
wait for Clk_period;
Addr <= "0001111000010";
Trees_din <= "00000011000000000101000100000100";
wait for Clk_period;
Addr <= "0001111000011";
Trees_din <= "00000000001001100001000011010101";
wait for Clk_period;
Addr <= "0001111000100";
Trees_din <= "00000000000100010001000011010101";
wait for Clk_period;
Addr <= "0001111000101";
Trees_din <= "00000000000000000001100100000100";
wait for Clk_period;
Addr <= "0001111000110";
Trees_din <= "00000000000111010001000011010101";
wait for Clk_period;
Addr <= "0001111000111";
Trees_din <= "00000000000011100001000011010101";
wait for Clk_period;
Addr <= "0001111001000";
Trees_din <= "00000111000000000100000100010000";
wait for Clk_period;
Addr <= "0001111001001";
Trees_din <= "00000100000000000100110100001000";
wait for Clk_period;
Addr <= "0001111001010";
Trees_din <= "00000100000000000000011000000100";
wait for Clk_period;
Addr <= "0001111001011";
Trees_din <= "00000000001100110001000011010101";
wait for Clk_period;
Addr <= "0001111001100";
Trees_din <= "00000000000011000001000011010101";
wait for Clk_period;
Addr <= "0001111001101";
Trees_din <= "00000011000000000110000100000100";
wait for Clk_period;
Addr <= "0001111001110";
Trees_din <= "00000000000000000001000011010101";
wait for Clk_period;
Addr <= "0001111001111";
Trees_din <= "00000000011000100001000011010101";
wait for Clk_period;
Addr <= "0001111010000";
Trees_din <= "00000010000000000010111100001000";
wait for Clk_period;
Addr <= "0001111010001";
Trees_din <= "00000011000000000000101100000100";
wait for Clk_period;
Addr <= "0001111010010";
Trees_din <= "00000000000111100001000011010101";
wait for Clk_period;
Addr <= "0001111010011";
Trees_din <= "00000000001111100001000011010101";
wait for Clk_period;
Addr <= "0001111010100";
Trees_din <= "00000010000000000001001100000100";
wait for Clk_period;
Addr <= "0001111010101";
Trees_din <= "00000000010001110001000011010101";
wait for Clk_period;
Addr <= "0001111010110";
Trees_din <= "00000000010101010001000011010101";
wait for Clk_period;
Addr <= "0001111010111";
Trees_din <= "00000001000000000001010000100000";
wait for Clk_period;
Addr <= "0001111011000";
Trees_din <= "00000010000000000110001000010000";
wait for Clk_period;
Addr <= "0001111011001";
Trees_din <= "00000111000000000100101100001000";
wait for Clk_period;
Addr <= "0001111011010";
Trees_din <= "00000000000000000000101000000100";
wait for Clk_period;
Addr <= "0001111011011";
Trees_din <= "00000000000011110001000011010101";
wait for Clk_period;
Addr <= "0001111011100";
Trees_din <= "00000000010001000001000011010101";
wait for Clk_period;
Addr <= "0001111011101";
Trees_din <= "00000111000000000110000100000100";
wait for Clk_period;
Addr <= "0001111011110";
Trees_din <= "00000000010011010001000011010101";
wait for Clk_period;
Addr <= "0001111011111";
Trees_din <= "00000000010000010001000011010101";
wait for Clk_period;
Addr <= "0001111100000";
Trees_din <= "00000010000000000001011100001000";
wait for Clk_period;
Addr <= "0001111100001";
Trees_din <= "00000101000000000001110100000100";
wait for Clk_period;
Addr <= "0001111100010";
Trees_din <= "00000000011001000001000011010101";
wait for Clk_period;
Addr <= "0001111100011";
Trees_din <= "00000000001011100001000011010101";
wait for Clk_period;
Addr <= "0001111100100";
Trees_din <= "00000111000000000011000000000100";
wait for Clk_period;
Addr <= "0001111100101";
Trees_din <= "00000000000100000001000011010101";
wait for Clk_period;
Addr <= "0001111100110";
Trees_din <= "00000000010010100001000011010101";
wait for Clk_period;
Addr <= "0001111100111";
Trees_din <= "00000011000000000011110000010000";
wait for Clk_period;
Addr <= "0001111101000";
Trees_din <= "00000001000000000100110000001000";
wait for Clk_period;
Addr <= "0001111101001";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "0001111101010";
Trees_din <= "00000000000111010001000011010101";
wait for Clk_period;
Addr <= "0001111101011";
Trees_din <= "00000000001110000001000011010101";
wait for Clk_period;
Addr <= "0001111101100";
Trees_din <= "00000111000000000101101000000100";
wait for Clk_period;
Addr <= "0001111101101";
Trees_din <= "00000000001000110001000011010101";
wait for Clk_period;
Addr <= "0001111101110";
Trees_din <= "00000000010001110001000011010101";
wait for Clk_period;
Addr <= "0001111101111";
Trees_din <= "00000101000000000000101100001000";
wait for Clk_period;
Addr <= "0001111110000";
Trees_din <= "00000001000000000011001100000100";
wait for Clk_period;
Addr <= "0001111110001";
Trees_din <= "00000000010110000001000011010101";
wait for Clk_period;
Addr <= "0001111110010";
Trees_din <= "00000000001100110001000011010101";
wait for Clk_period;
Addr <= "0001111110011";
Trees_din <= "00000100000000000010100000000100";
wait for Clk_period;
Addr <= "0001111110100";
Trees_din <= "00000000001111110001000011010101";
wait for Clk_period;
Addr <= "0001111110101";
Trees_din <= "00000000010101000001000011010101";
wait for Clk_period;
Addr <= "0001111110110";
Trees_din <= "00000111000000000010011101000000";
wait for Clk_period;
Addr <= "0001111110111";
Trees_din <= "00000101000000000100001000100000";
wait for Clk_period;
Addr <= "0001111111000";
Trees_din <= "00000110000000000100100100010000";
wait for Clk_period;
Addr <= "0001111111001";
Trees_din <= "00000100000000000010000000001000";
wait for Clk_period;
Addr <= "0001111111010";
Trees_din <= "00000011000000000011001000000100";
wait for Clk_period;
Addr <= "0001111111011";
Trees_din <= "00000000001000010001000011010101";
wait for Clk_period;
Addr <= "0001111111100";
Trees_din <= "00000000001011000001000011010101";
wait for Clk_period;
Addr <= "0001111111101";
Trees_din <= "00000000000000000000010100000100";
wait for Clk_period;
Addr <= "0001111111110";
Trees_din <= "00000000001111100001000011010101";
wait for Clk_period;
Addr <= "0001111111111";
Trees_din <= "00000000000000000001000011010101";
wait for Clk_period;
Addr <= "0010000000000";
Trees_din <= "00000111000000000101110100001000";
wait for Clk_period;
Addr <= "0010000000001";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "0010000000010";
Trees_din <= "00000000010000100001000011010101";
wait for Clk_period;
Addr <= "0010000000011";
Trees_din <= "00000000001001110001000011010101";
wait for Clk_period;
Addr <= "0010000000100";
Trees_din <= "00000101000000000010011100000100";
wait for Clk_period;
Addr <= "0010000000101";
Trees_din <= "00000000010101010001000011010101";
wait for Clk_period;
Addr <= "0010000000110";
Trees_din <= "00000000000000100001000011010101";
wait for Clk_period;
Addr <= "0010000000111";
Trees_din <= "00000011000000000000001100010000";
wait for Clk_period;
Addr <= "0010000001000";
Trees_din <= "00000011000000000001011000001000";
wait for Clk_period;
Addr <= "0010000001001";
Trees_din <= "00000110000000000000011100000100";
wait for Clk_period;
Addr <= "0010000001010";
Trees_din <= "00000000001101100001000011010101";
wait for Clk_period;
Addr <= "0010000001011";
Trees_din <= "00000000000100000001000011010101";
wait for Clk_period;
Addr <= "0010000001100";
Trees_din <= "00000101000000000010101100000100";
wait for Clk_period;
Addr <= "0010000001101";
Trees_din <= "00000000000111100001000011010101";
wait for Clk_period;
Addr <= "0010000001110";
Trees_din <= "00000000000100100001000011010101";
wait for Clk_period;
Addr <= "0010000001111";
Trees_din <= "00000110000000000101111100001000";
wait for Clk_period;
Addr <= "0010000010000";
Trees_din <= "00000001000000000011010000000100";
wait for Clk_period;
Addr <= "0010000010001";
Trees_din <= "00000000011001000001000011010101";
wait for Clk_period;
Addr <= "0010000010010";
Trees_din <= "00000000010000010001000011010101";
wait for Clk_period;
Addr <= "0010000010011";
Trees_din <= "00000111000000000000111000000100";
wait for Clk_period;
Addr <= "0010000010100";
Trees_din <= "00000000001111000001000011010101";
wait for Clk_period;
Addr <= "0010000010101";
Trees_din <= "00000000000011010001000011010101";
wait for Clk_period;
Addr <= "0010000010110";
Trees_din <= "00000010000000000000101000100000";
wait for Clk_period;
Addr <= "0010000010111";
Trees_din <= "00000100000000000110000100010000";
wait for Clk_period;
Addr <= "0010000011000";
Trees_din <= "00000001000000000110010000001000";
wait for Clk_period;
Addr <= "0010000011001";
Trees_din <= "00000100000000000010100000000100";
wait for Clk_period;
Addr <= "0010000011010";
Trees_din <= "00000000001001010001000011010101";
wait for Clk_period;
Addr <= "0010000011011";
Trees_din <= "00000000000000000001000011010101";
wait for Clk_period;
Addr <= "0010000011100";
Trees_din <= "00000001000000000101010100000100";
wait for Clk_period;
Addr <= "0010000011101";
Trees_din <= "00000000010001110001000011010101";
wait for Clk_period;
Addr <= "0010000011110";
Trees_din <= "00000000010010000001000011010101";
wait for Clk_period;
Addr <= "0010000011111";
Trees_din <= "00000101000000000001110100001000";
wait for Clk_period;
Addr <= "0010000100000";
Trees_din <= "00000000000000000011001000000100";
wait for Clk_period;
Addr <= "0010000100001";
Trees_din <= "00000000010101110001000011010101";
wait for Clk_period;
Addr <= "0010000100010";
Trees_din <= "00000000000000000001000011010101";
wait for Clk_period;
Addr <= "0010000100011";
Trees_din <= "00000011000000000100100100000100";
wait for Clk_period;
Addr <= "0010000100100";
Trees_din <= "00000000000111110001000011010101";
wait for Clk_period;
Addr <= "0010000100101";
Trees_din <= "00000000011000000001000011010101";
wait for Clk_period;
Addr <= "0010000100110";
Trees_din <= "00000000000000000001001000010000";
wait for Clk_period;
Addr <= "0010000100111";
Trees_din <= "00000011000000000011111000001000";
wait for Clk_period;
Addr <= "0010000101000";
Trees_din <= "00000011000000000100110100000100";
wait for Clk_period;
Addr <= "0010000101001";
Trees_din <= "00000000001100110001000011010101";
wait for Clk_period;
Addr <= "0010000101010";
Trees_din <= "00000000000011010001000011010101";
wait for Clk_period;
Addr <= "0010000101011";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "0010000101100";
Trees_din <= "00000000010101100001000011010101";
wait for Clk_period;
Addr <= "0010000101101";
Trees_din <= "00000000001101110001000011010101";
wait for Clk_period;
Addr <= "0010000101110";
Trees_din <= "00000000000000000100011100001000";
wait for Clk_period;
Addr <= "0010000101111";
Trees_din <= "00000111000000000100110100000100";
wait for Clk_period;
Addr <= "0010000110000";
Trees_din <= "00000000001101000001000011010101";
wait for Clk_period;
Addr <= "0010000110001";
Trees_din <= "00000000011000100001000011010101";
wait for Clk_period;
Addr <= "0010000110010";
Trees_din <= "00000101000000000100010000000100";
wait for Clk_period;
Addr <= "0010000110011";
Trees_din <= "00000000010001110001000011010101";
wait for Clk_period;
Addr <= "0010000110100";
Trees_din <= "00000000010010010001000011010101";
wait for Clk_period;



----------tree 8-------------------

Addr <= "0010000110101";
Trees_din <= "00000101000000000100111110000000";
wait for Clk_period;
Addr <= "0010000110110";
Trees_din <= "00000111000000000100100001000000";
wait for Clk_period;
Addr <= "0010000110111";
Trees_din <= "00000010000000000010110000100000";
wait for Clk_period;
Addr <= "0010000111000";
Trees_din <= "00000110000000000100110000010000";
wait for Clk_period;
Addr <= "0010000111001";
Trees_din <= "00000011000000000101010100001000";
wait for Clk_period;
Addr <= "0010000111010";
Trees_din <= "00000101000000000110010000000100";
wait for Clk_period;
Addr <= "0010000111011";
Trees_din <= "00000000010111000001001011010001";
wait for Clk_period;
Addr <= "0010000111100";
Trees_din <= "00000000001100110001001011010001";
wait for Clk_period;
Addr <= "0010000111101";
Trees_din <= "00000101000000000010010100000100";
wait for Clk_period;
Addr <= "0010000111110";
Trees_din <= "00000000001010000001001011010001";
wait for Clk_period;
Addr <= "0010000111111";
Trees_din <= "00000000010010100001001011010001";
wait for Clk_period;
Addr <= "0010001000000";
Trees_din <= "00000111000000000101001100001000";
wait for Clk_period;
Addr <= "0010001000001";
Trees_din <= "00000010000000000000101000000100";
wait for Clk_period;
Addr <= "0010001000010";
Trees_din <= "00000000001000000001001011010001";
wait for Clk_period;
Addr <= "0010001000011";
Trees_din <= "00000000000000100001001011010001";
wait for Clk_period;
Addr <= "0010001000100";
Trees_din <= "00000100000000000001001100000100";
wait for Clk_period;
Addr <= "0010001000101";
Trees_din <= "00000000010111010001001011010001";
wait for Clk_period;
Addr <= "0010001000110";
Trees_din <= "00000000000100110001001011010001";
wait for Clk_period;
Addr <= "0010001000111";
Trees_din <= "00000100000000000010001000010000";
wait for Clk_period;
Addr <= "0010001001000";
Trees_din <= "00000110000000000001011100001000";
wait for Clk_period;
Addr <= "0010001001001";
Trees_din <= "00000001000000000000110100000100";
wait for Clk_period;
Addr <= "0010001001010";
Trees_din <= "00000000010101010001001011010001";
wait for Clk_period;
Addr <= "0010001001011";
Trees_din <= "00000000000100100001001011010001";
wait for Clk_period;
Addr <= "0010001001100";
Trees_din <= "00000010000000000000110100000100";
wait for Clk_period;
Addr <= "0010001001101";
Trees_din <= "00000000001110000001001011010001";
wait for Clk_period;
Addr <= "0010001001110";
Trees_din <= "00000000000010010001001011010001";
wait for Clk_period;
Addr <= "0010001001111";
Trees_din <= "00000111000000000000011100001000";
wait for Clk_period;
Addr <= "0010001010000";
Trees_din <= "00000100000000000110001000000100";
wait for Clk_period;
Addr <= "0010001010001";
Trees_din <= "00000000001010010001001011010001";
wait for Clk_period;
Addr <= "0010001010010";
Trees_din <= "00000000001110110001001011010001";
wait for Clk_period;
Addr <= "0010001010011";
Trees_din <= "00000001000000000100101000000100";
wait for Clk_period;
Addr <= "0010001010100";
Trees_din <= "00000000000010100001001011010001";
wait for Clk_period;
Addr <= "0010001010101";
Trees_din <= "00000000000100000001001011010001";
wait for Clk_period;
Addr <= "0010001010110";
Trees_din <= "00000010000000000001111100100000";
wait for Clk_period;
Addr <= "0010001010111";
Trees_din <= "00000100000000000000110100010000";
wait for Clk_period;
Addr <= "0010001011000";
Trees_din <= "00000110000000000100111100001000";
wait for Clk_period;
Addr <= "0010001011001";
Trees_din <= "00000010000000000100110000000100";
wait for Clk_period;
Addr <= "0010001011010";
Trees_din <= "00000000001100110001001011010001";
wait for Clk_period;
Addr <= "0010001011011";
Trees_din <= "00000000001000100001001011010001";
wait for Clk_period;
Addr <= "0010001011100";
Trees_din <= "00000011000000000000111000000100";
wait for Clk_period;
Addr <= "0010001011101";
Trees_din <= "00000000001001100001001011010001";
wait for Clk_period;
Addr <= "0010001011110";
Trees_din <= "00000000001110000001001011010001";
wait for Clk_period;
Addr <= "0010001011111";
Trees_din <= "00000010000000000100011000001000";
wait for Clk_period;
Addr <= "0010001100000";
Trees_din <= "00000000000000000011001100000100";
wait for Clk_period;
Addr <= "0010001100001";
Trees_din <= "00000000001001100001001011010001";
wait for Clk_period;
Addr <= "0010001100010";
Trees_din <= "00000000001010010001001011010001";
wait for Clk_period;
Addr <= "0010001100011";
Trees_din <= "00000010000000000101110100000100";
wait for Clk_period;
Addr <= "0010001100100";
Trees_din <= "00000000001111010001001011010001";
wait for Clk_period;
Addr <= "0010001100101";
Trees_din <= "00000000011000010001001011010001";
wait for Clk_period;
Addr <= "0010001100110";
Trees_din <= "00000001000000000010111100010000";
wait for Clk_period;
Addr <= "0010001100111";
Trees_din <= "00000101000000000011101000001000";
wait for Clk_period;
Addr <= "0010001101000";
Trees_din <= "00000100000000000011011100000100";
wait for Clk_period;
Addr <= "0010001101001";
Trees_din <= "00000000010101100001001011010001";
wait for Clk_period;
Addr <= "0010001101010";
Trees_din <= "00000000001100000001001011010001";
wait for Clk_period;
Addr <= "0010001101011";
Trees_din <= "00000011000000000000011000000100";
wait for Clk_period;
Addr <= "0010001101100";
Trees_din <= "00000000000000010001001011010001";
wait for Clk_period;
Addr <= "0010001101101";
Trees_din <= "00000000010100000001001011010001";
wait for Clk_period;
Addr <= "0010001101110";
Trees_din <= "00000110000000000001101000001000";
wait for Clk_period;
Addr <= "0010001101111";
Trees_din <= "00000111000000000011100100000100";
wait for Clk_period;
Addr <= "0010001110000";
Trees_din <= "00000000000100010001001011010001";
wait for Clk_period;
Addr <= "0010001110001";
Trees_din <= "00000000001001100001001011010001";
wait for Clk_period;
Addr <= "0010001110010";
Trees_din <= "00000001000000000101111000000100";
wait for Clk_period;
Addr <= "0010001110011";
Trees_din <= "00000000000111100001001011010001";
wait for Clk_period;
Addr <= "0010001110100";
Trees_din <= "00000000010111110001001011010001";
wait for Clk_period;
Addr <= "0010001110101";
Trees_din <= "00000100000000000100100101000000";
wait for Clk_period;
Addr <= "0010001110110";
Trees_din <= "00000000000000000101010000100000";
wait for Clk_period;
Addr <= "0010001110111";
Trees_din <= "00000010000000000110001000010000";
wait for Clk_period;
Addr <= "0010001111000";
Trees_din <= "00000001000000000001100000001000";
wait for Clk_period;
Addr <= "0010001111001";
Trees_din <= "00000010000000000010110100000100";
wait for Clk_period;
Addr <= "0010001111010";
Trees_din <= "00000000000001100001001011010001";
wait for Clk_period;
Addr <= "0010001111011";
Trees_din <= "00000000000101110001001011010001";
wait for Clk_period;
Addr <= "0010001111100";
Trees_din <= "00000011000000000000011000000100";
wait for Clk_period;
Addr <= "0010001111101";
Trees_din <= "00000000010000110001001011010001";
wait for Clk_period;
Addr <= "0010001111110";
Trees_din <= "00000000000011000001001011010001";
wait for Clk_period;
Addr <= "0010001111111";
Trees_din <= "00000011000000000000101000001000";
wait for Clk_period;
Addr <= "0010010000000";
Trees_din <= "00000111000000000101000000000100";
wait for Clk_period;
Addr <= "0010010000001";
Trees_din <= "00000000001110010001001011010001";
wait for Clk_period;
Addr <= "0010010000010";
Trees_din <= "00000000010001110001001011010001";
wait for Clk_period;
Addr <= "0010010000011";
Trees_din <= "00000000000000000000110000000100";
wait for Clk_period;
Addr <= "0010010000100";
Trees_din <= "00000000000101110001001011010001";
wait for Clk_period;
Addr <= "0010010000101";
Trees_din <= "00000000010111000001001011010001";
wait for Clk_period;
Addr <= "0010010000110";
Trees_din <= "00000000000000000100000000010000";
wait for Clk_period;
Addr <= "0010010000111";
Trees_din <= "00000111000000000100010000001000";
wait for Clk_period;
Addr <= "0010010001000";
Trees_din <= "00000011000000000000110000000100";
wait for Clk_period;
Addr <= "0010010001001";
Trees_din <= "00000000001001110001001011010001";
wait for Clk_period;
Addr <= "0010010001010";
Trees_din <= "00000000000110110001001011010001";
wait for Clk_period;
Addr <= "0010010001011";
Trees_din <= "00000101000000000011000100000100";
wait for Clk_period;
Addr <= "0010010001100";
Trees_din <= "00000000000111010001001011010001";
wait for Clk_period;
Addr <= "0010010001101";
Trees_din <= "00000000010111110001001011010001";
wait for Clk_period;
Addr <= "0010010001110";
Trees_din <= "00000110000000000101100000001000";
wait for Clk_period;
Addr <= "0010010001111";
Trees_din <= "00000001000000000010010000000100";
wait for Clk_period;
Addr <= "0010010010000";
Trees_din <= "00000000001111100001001011010001";
wait for Clk_period;
Addr <= "0010010010001";
Trees_din <= "00000000001110100001001011010001";
wait for Clk_period;
Addr <= "0010010010010";
Trees_din <= "00000111000000000001010000000100";
wait for Clk_period;
Addr <= "0010010010011";
Trees_din <= "00000000001100010001001011010001";
wait for Clk_period;
Addr <= "0010010010100";
Trees_din <= "00000000001111000001001011010001";
wait for Clk_period;
Addr <= "0010010010101";
Trees_din <= "00000100000000000011000100100000";
wait for Clk_period;
Addr <= "0010010010110";
Trees_din <= "00000111000000000011100100010000";
wait for Clk_period;
Addr <= "0010010010111";
Trees_din <= "00000011000000000001001100001000";
wait for Clk_period;
Addr <= "0010010011000";
Trees_din <= "00000010000000000101110100000100";
wait for Clk_period;
Addr <= "0010010011001";
Trees_din <= "00000000000111000001001011010001";
wait for Clk_period;
Addr <= "0010010011010";
Trees_din <= "00000000010111100001001011010001";
wait for Clk_period;
Addr <= "0010010011011";
Trees_din <= "00000000000000000010111100000100";
wait for Clk_period;
Addr <= "0010010011100";
Trees_din <= "00000000010010100001001011010001";
wait for Clk_period;
Addr <= "0010010011101";
Trees_din <= "00000000000011000001001011010001";
wait for Clk_period;
Addr <= "0010010011110";
Trees_din <= "00000110000000000100010000001000";
wait for Clk_period;
Addr <= "0010010011111";
Trees_din <= "00000111000000000101100100000100";
wait for Clk_period;
Addr <= "0010010100000";
Trees_din <= "00000000000111110001001011010001";
wait for Clk_period;
Addr <= "0010010100001";
Trees_din <= "00000000000100010001001011010001";
wait for Clk_period;
Addr <= "0010010100010";
Trees_din <= "00000101000000000001110100000100";
wait for Clk_period;
Addr <= "0010010100011";
Trees_din <= "00000000011000110001001011010001";
wait for Clk_period;
Addr <= "0010010100100";
Trees_din <= "00000000010110100001001011010001";
wait for Clk_period;
Addr <= "0010010100101";
Trees_din <= "00000000000000000001101000010000";
wait for Clk_period;
Addr <= "0010010100110";
Trees_din <= "00000011000000000011110000001000";
wait for Clk_period;
Addr <= "0010010100111";
Trees_din <= "00000000000000000000010100000100";
wait for Clk_period;
Addr <= "0010010101000";
Trees_din <= "00000000010110010001001011010001";
wait for Clk_period;
Addr <= "0010010101001";
Trees_din <= "00000000001100100001001011010001";
wait for Clk_period;
Addr <= "0010010101010";
Trees_din <= "00000000000000000100110000000100";
wait for Clk_period;
Addr <= "0010010101011";
Trees_din <= "00000000000000110001001011010001";
wait for Clk_period;
Addr <= "0010010101100";
Trees_din <= "00000000010010110001001011010001";
wait for Clk_period;
Addr <= "0010010101101";
Trees_din <= "00000011000000000000111000001000";
wait for Clk_period;
Addr <= "0010010101110";
Trees_din <= "00000110000000000001011100000100";
wait for Clk_period;
Addr <= "0010010101111";
Trees_din <= "00000000010001100001001011010001";
wait for Clk_period;
Addr <= "0010010110000";
Trees_din <= "00000000000101010001001011010001";
wait for Clk_period;
Addr <= "0010010110001";
Trees_din <= "00000011000000000000001100000100";
wait for Clk_period;
Addr <= "0010010110010";
Trees_din <= "00000000010010110001001011010001";
wait for Clk_period;
Addr <= "0010010110011";
Trees_din <= "00000000010110000001001011010001";
wait for Clk_period;



----------tree 9-------------------

Addr <= "0010010110100";
Trees_din <= "00000001000000000001110010000000";
wait for Clk_period;
Addr <= "0010010110101";
Trees_din <= "00000011000000000010001001000000";
wait for Clk_period;
Addr <= "0010010110110";
Trees_din <= "00000101000000000010110100100000";
wait for Clk_period;
Addr <= "0010010110111";
Trees_din <= "00000000000000000011100000010000";
wait for Clk_period;
Addr <= "0010010111000";
Trees_din <= "00000010000000000110001100001000";
wait for Clk_period;
Addr <= "0010010111001";
Trees_din <= "00000110000000000011001100000100";
wait for Clk_period;
Addr <= "0010010111010";
Trees_din <= "00000000000010000001010011001101";
wait for Clk_period;
Addr <= "0010010111011";
Trees_din <= "00000000001110110001010011001101";
wait for Clk_period;
Addr <= "0010010111100";
Trees_din <= "00000001000000000010101100000100";
wait for Clk_period;
Addr <= "0010010111101";
Trees_din <= "00000000000110000001010011001101";
wait for Clk_period;
Addr <= "0010010111110";
Trees_din <= "00000000010111100001010011001101";
wait for Clk_period;
Addr <= "0010010111111";
Trees_din <= "00000001000000000000010000001000";
wait for Clk_period;
Addr <= "0010011000000";
Trees_din <= "00000001000000000000101100000100";
wait for Clk_period;
Addr <= "0010011000001";
Trees_din <= "00000000001101110001010011001101";
wait for Clk_period;
Addr <= "0010011000010";
Trees_din <= "00000000010000000001010011001101";
wait for Clk_period;
Addr <= "0010011000011";
Trees_din <= "00000001000000000001101000000100";
wait for Clk_period;
Addr <= "0010011000100";
Trees_din <= "00000000001001000001010011001101";
wait for Clk_period;
Addr <= "0010011000101";
Trees_din <= "00000000010110110001010011001101";
wait for Clk_period;
Addr <= "0010011000110";
Trees_din <= "00000111000000000100011000010000";
wait for Clk_period;
Addr <= "0010011000111";
Trees_din <= "00000100000000000100111100001000";
wait for Clk_period;
Addr <= "0010011001000";
Trees_din <= "00000111000000000000011100000100";
wait for Clk_period;
Addr <= "0010011001001";
Trees_din <= "00000000000100110001010011001101";
wait for Clk_period;
Addr <= "0010011001010";
Trees_din <= "00000000000111100001010011001101";
wait for Clk_period;
Addr <= "0010011001011";
Trees_din <= "00000001000000000001010000000100";
wait for Clk_period;
Addr <= "0010011001100";
Trees_din <= "00000000010110010001010011001101";
wait for Clk_period;
Addr <= "0010011001101";
Trees_din <= "00000000000001110001010011001101";
wait for Clk_period;
Addr <= "0010011001110";
Trees_din <= "00000011000000000101000100001000";
wait for Clk_period;
Addr <= "0010011001111";
Trees_din <= "00000010000000000110000000000100";
wait for Clk_period;
Addr <= "0010011010000";
Trees_din <= "00000000001010010001010011001101";
wait for Clk_period;
Addr <= "0010011010001";
Trees_din <= "00000000001001010001010011001101";
wait for Clk_period;
Addr <= "0010011010010";
Trees_din <= "00000111000000000000001000000100";
wait for Clk_period;
Addr <= "0010011010011";
Trees_din <= "00000000010100000001010011001101";
wait for Clk_period;
Addr <= "0010011010100";
Trees_din <= "00000000010010010001010011001101";
wait for Clk_period;
Addr <= "0010011010101";
Trees_din <= "00000100000000000100001100100000";
wait for Clk_period;
Addr <= "0010011010110";
Trees_din <= "00000101000000000011001000010000";
wait for Clk_period;
Addr <= "0010011010111";
Trees_din <= "00000000000000000000101100001000";
wait for Clk_period;
Addr <= "0010011011000";
Trees_din <= "00000011000000000000001000000100";
wait for Clk_period;
Addr <= "0010011011001";
Trees_din <= "00000000000101010001010011001101";
wait for Clk_period;
Addr <= "0010011011010";
Trees_din <= "00000000000110100001010011001101";
wait for Clk_period;
Addr <= "0010011011011";
Trees_din <= "00000010000000000010000000000100";
wait for Clk_period;
Addr <= "0010011011100";
Trees_din <= "00000000010011010001010011001101";
wait for Clk_period;
Addr <= "0010011011101";
Trees_din <= "00000000000001110001010011001101";
wait for Clk_period;
Addr <= "0010011011110";
Trees_din <= "00000010000000000000111100001000";
wait for Clk_period;
Addr <= "0010011011111";
Trees_din <= "00000001000000000001001000000100";
wait for Clk_period;
Addr <= "0010011100000";
Trees_din <= "00000000000110000001010011001101";
wait for Clk_period;
Addr <= "0010011100001";
Trees_din <= "00000000000111000001010011001101";
wait for Clk_period;
Addr <= "0010011100010";
Trees_din <= "00000111000000000001101100000100";
wait for Clk_period;
Addr <= "0010011100011";
Trees_din <= "00000000000100010001010011001101";
wait for Clk_period;
Addr <= "0010011100100";
Trees_din <= "00000000000001110001010011001101";
wait for Clk_period;
Addr <= "0010011100101";
Trees_din <= "00000101000000000110001000010000";
wait for Clk_period;
Addr <= "0010011100110";
Trees_din <= "00000011000000000101110000001000";
wait for Clk_period;
Addr <= "0010011100111";
Trees_din <= "00000000000000000101001000000100";
wait for Clk_period;
Addr <= "0010011101000";
Trees_din <= "00000000011000000001010011001101";
wait for Clk_period;
Addr <= "0010011101001";
Trees_din <= "00000000010101100001010011001101";
wait for Clk_period;
Addr <= "0010011101010";
Trees_din <= "00000101000000000011000100000100";
wait for Clk_period;
Addr <= "0010011101011";
Trees_din <= "00000000000010010001010011001101";
wait for Clk_period;
Addr <= "0010011101100";
Trees_din <= "00000000000101110001010011001101";
wait for Clk_period;
Addr <= "0010011101101";
Trees_din <= "00000011000000000110010000001000";
wait for Clk_period;
Addr <= "0010011101110";
Trees_din <= "00000111000000000001011100000100";
wait for Clk_period;
Addr <= "0010011101111";
Trees_din <= "00000000010110110001010011001101";
wait for Clk_period;
Addr <= "0010011110000";
Trees_din <= "00000000000000100001010011001101";
wait for Clk_period;
Addr <= "0010011110001";
Trees_din <= "00000110000000000001011100000100";
wait for Clk_period;
Addr <= "0010011110010";
Trees_din <= "00000000010100010001010011001101";
wait for Clk_period;
Addr <= "0010011110011";
Trees_din <= "00000000000101100001010011001101";
wait for Clk_period;
Addr <= "0010011110100";
Trees_din <= "00000110000000000100001101000000";
wait for Clk_period;
Addr <= "0010011110101";
Trees_din <= "00000100000000000001100000100000";
wait for Clk_period;
Addr <= "0010011110110";
Trees_din <= "00000010000000000000111100010000";
wait for Clk_period;
Addr <= "0010011110111";
Trees_din <= "00000110000000000101001000001000";
wait for Clk_period;
Addr <= "0010011111000";
Trees_din <= "00000001000000000101101000000100";
wait for Clk_period;
Addr <= "0010011111001";
Trees_din <= "00000000001001100001010011001101";
wait for Clk_period;
Addr <= "0010011111010";
Trees_din <= "00000000000111010001010011001101";
wait for Clk_period;
Addr <= "0010011111011";
Trees_din <= "00000100000000000110001000000100";
wait for Clk_period;
Addr <= "0010011111100";
Trees_din <= "00000000010100000001010011001101";
wait for Clk_period;
Addr <= "0010011111101";
Trees_din <= "00000000000100000001010011001101";
wait for Clk_period;
Addr <= "0010011111110";
Trees_din <= "00000010000000000010011100001000";
wait for Clk_period;
Addr <= "0010011111111";
Trees_din <= "00000001000000000001100000000100";
wait for Clk_period;
Addr <= "0010100000000";
Trees_din <= "00000000000011000001010011001101";
wait for Clk_period;
Addr <= "0010100000001";
Trees_din <= "00000000010000110001010011001101";
wait for Clk_period;
Addr <= "0010100000010";
Trees_din <= "00000000000000000000111000000100";
wait for Clk_period;
Addr <= "0010100000011";
Trees_din <= "00000000010111100001010011001101";
wait for Clk_period;
Addr <= "0010100000100";
Trees_din <= "00000000010001000001010011001101";
wait for Clk_period;
Addr <= "0010100000101";
Trees_din <= "00000110000000000001001000010000";
wait for Clk_period;
Addr <= "0010100000110";
Trees_din <= "00000000000000000101100000001000";
wait for Clk_period;
Addr <= "0010100000111";
Trees_din <= "00000011000000000100001000000100";
wait for Clk_period;
Addr <= "0010100001000";
Trees_din <= "00000000000010110001010011001101";
wait for Clk_period;
Addr <= "0010100001001";
Trees_din <= "00000000000011000001010011001101";
wait for Clk_period;
Addr <= "0010100001010";
Trees_din <= "00000101000000000001111000000100";
wait for Clk_period;
Addr <= "0010100001011";
Trees_din <= "00000000010010110001010011001101";
wait for Clk_period;
Addr <= "0010100001100";
Trees_din <= "00000000000100010001010011001101";
wait for Clk_period;
Addr <= "0010100001101";
Trees_din <= "00000000000000000010011100001000";
wait for Clk_period;
Addr <= "0010100001110";
Trees_din <= "00000110000000000010101000000100";
wait for Clk_period;
Addr <= "0010100001111";
Trees_din <= "00000000010111100001010011001101";
wait for Clk_period;
Addr <= "0010100010000";
Trees_din <= "00000000010011010001010011001101";
wait for Clk_period;
Addr <= "0010100010001";
Trees_din <= "00000101000000000010110000000100";
wait for Clk_period;
Addr <= "0010100010010";
Trees_din <= "00000000010110100001010011001101";
wait for Clk_period;
Addr <= "0010100010011";
Trees_din <= "00000000000000010001010011001101";
wait for Clk_period;
Addr <= "0010100010100";
Trees_din <= "00000101000000000001000000100000";
wait for Clk_period;
Addr <= "0010100010101";
Trees_din <= "00000100000000000100010100010000";
wait for Clk_period;
Addr <= "0010100010110";
Trees_din <= "00000100000000000100010000001000";
wait for Clk_period;
Addr <= "0010100010111";
Trees_din <= "00000010000000000011111100000100";
wait for Clk_period;
Addr <= "0010100011000";
Trees_din <= "00000000001100000001010011001101";
wait for Clk_period;
Addr <= "0010100011001";
Trees_din <= "00000000010101100001010011001101";
wait for Clk_period;
Addr <= "0010100011010";
Trees_din <= "00000001000000000011010100000100";
wait for Clk_period;
Addr <= "0010100011011";
Trees_din <= "00000000001011000001010011001101";
wait for Clk_period;
Addr <= "0010100011100";
Trees_din <= "00000000001011100001010011001101";
wait for Clk_period;
Addr <= "0010100011101";
Trees_din <= "00000011000000000000110100001000";
wait for Clk_period;
Addr <= "0010100011110";
Trees_din <= "00000111000000000101100000000100";
wait for Clk_period;
Addr <= "0010100011111";
Trees_din <= "00000000000001110001010011001101";
wait for Clk_period;
Addr <= "0010100100000";
Trees_din <= "00000000000101100001010011001101";
wait for Clk_period;
Addr <= "0010100100001";
Trees_din <= "00000000000000000001110100000100";
wait for Clk_period;
Addr <= "0010100100010";
Trees_din <= "00000000010111010001010011001101";
wait for Clk_period;
Addr <= "0010100100011";
Trees_din <= "00000000000010000001010011001101";
wait for Clk_period;
Addr <= "0010100100100";
Trees_din <= "00000110000000000011011000010000";
wait for Clk_period;
Addr <= "0010100100101";
Trees_din <= "00000010000000000000000100001000";
wait for Clk_period;
Addr <= "0010100100110";
Trees_din <= "00000111000000000101100000000100";
wait for Clk_period;
Addr <= "0010100100111";
Trees_din <= "00000000001011000001010011001101";
wait for Clk_period;
Addr <= "0010100101000";
Trees_din <= "00000000010111110001010011001101";
wait for Clk_period;
Addr <= "0010100101001";
Trees_din <= "00000001000000000000001000000100";
wait for Clk_period;
Addr <= "0010100101010";
Trees_din <= "00000000000001010001010011001101";
wait for Clk_period;
Addr <= "0010100101011";
Trees_din <= "00000000010011100001010011001101";
wait for Clk_period;
Addr <= "0010100101100";
Trees_din <= "00000011000000000011111100001000";
wait for Clk_period;
Addr <= "0010100101101";
Trees_din <= "00000001000000000101111100000100";
wait for Clk_period;
Addr <= "0010100101110";
Trees_din <= "00000000010000100001010011001101";
wait for Clk_period;
Addr <= "0010100101111";
Trees_din <= "00000000010111000001010011001101";
wait for Clk_period;
Addr <= "0010100110000";
Trees_din <= "00000011000000000011000000000100";
wait for Clk_period;
Addr <= "0010100110001";
Trees_din <= "00000000010000100001010011001101";
wait for Clk_period;
Addr <= "0010100110010";
Trees_din <= "00000000000101000001010011001101";
wait for Clk_period;



----------tree 10-------------------

Addr <= "0010100110011";
Trees_din <= "00000000000000000010111110000000";
wait for Clk_period;
Addr <= "0010100110100";
Trees_din <= "00000000000000000011010001000000";
wait for Clk_period;
Addr <= "0010100110101";
Trees_din <= "00000101000000000001110000100000";
wait for Clk_period;
Addr <= "0010100110110";
Trees_din <= "00000101000000000101111100010000";
wait for Clk_period;
Addr <= "0010100110111";
Trees_din <= "00000001000000000110000100001000";
wait for Clk_period;
Addr <= "0010100111000";
Trees_din <= "00000001000000000001000100000100";
wait for Clk_period;
Addr <= "0010100111001";
Trees_din <= "00000000001000000001011011001001";
wait for Clk_period;
Addr <= "0010100111010";
Trees_din <= "00000000000110000001011011001001";
wait for Clk_period;
Addr <= "0010100111011";
Trees_din <= "00000100000000000011110100000100";
wait for Clk_period;
Addr <= "0010100111100";
Trees_din <= "00000000000101010001011011001001";
wait for Clk_period;
Addr <= "0010100111101";
Trees_din <= "00000000001111010001011011001001";
wait for Clk_period;
Addr <= "0010100111110";
Trees_din <= "00000010000000000100010100001000";
wait for Clk_period;
Addr <= "0010100111111";
Trees_din <= "00000010000000000100010100000100";
wait for Clk_period;
Addr <= "0010101000000";
Trees_din <= "00000000010000110001011011001001";
wait for Clk_period;
Addr <= "0010101000001";
Trees_din <= "00000000001000110001011011001001";
wait for Clk_period;
Addr <= "0010101000010";
Trees_din <= "00000001000000000101010000000100";
wait for Clk_period;
Addr <= "0010101000011";
Trees_din <= "00000000010001000001011011001001";
wait for Clk_period;
Addr <= "0010101000100";
Trees_din <= "00000000010010100001011011001001";
wait for Clk_period;
Addr <= "0010101000101";
Trees_din <= "00000111000000000101111100010000";
wait for Clk_period;
Addr <= "0010101000110";
Trees_din <= "00000010000000000010100100001000";
wait for Clk_period;
Addr <= "0010101000111";
Trees_din <= "00000010000000000011111000000100";
wait for Clk_period;
Addr <= "0010101001000";
Trees_din <= "00000000000001100001011011001001";
wait for Clk_period;
Addr <= "0010101001001";
Trees_din <= "00000000010001110001011011001001";
wait for Clk_period;
Addr <= "0010101001010";
Trees_din <= "00000100000000000011101100000100";
wait for Clk_period;
Addr <= "0010101001011";
Trees_din <= "00000000000010110001011011001001";
wait for Clk_period;
Addr <= "0010101001100";
Trees_din <= "00000000001110010001011011001001";
wait for Clk_period;
Addr <= "0010101001101";
Trees_din <= "00000011000000000010110000001000";
wait for Clk_period;
Addr <= "0010101001110";
Trees_din <= "00000010000000000010110000000100";
wait for Clk_period;
Addr <= "0010101001111";
Trees_din <= "00000000010011100001011011001001";
wait for Clk_period;
Addr <= "0010101010000";
Trees_din <= "00000000000111110001011011001001";
wait for Clk_period;
Addr <= "0010101010001";
Trees_din <= "00000100000000000100010100000100";
wait for Clk_period;
Addr <= "0010101010010";
Trees_din <= "00000000010000000001011011001001";
wait for Clk_period;
Addr <= "0010101010011";
Trees_din <= "00000000001011110001011011001001";
wait for Clk_period;
Addr <= "0010101010100";
Trees_din <= "00000101000000000100000100100000";
wait for Clk_period;
Addr <= "0010101010101";
Trees_din <= "00000111000000000000000000010000";
wait for Clk_period;
Addr <= "0010101010110";
Trees_din <= "00000001000000000011000000001000";
wait for Clk_period;
Addr <= "0010101010111";
Trees_din <= "00000111000000000001000100000100";
wait for Clk_period;
Addr <= "0010101011000";
Trees_din <= "00000000001001100001011011001001";
wait for Clk_period;
Addr <= "0010101011001";
Trees_din <= "00000000001001000001011011001001";
wait for Clk_period;
Addr <= "0010101011010";
Trees_din <= "00000001000000000110010000000100";
wait for Clk_period;
Addr <= "0010101011011";
Trees_din <= "00000000001111100001011011001001";
wait for Clk_period;
Addr <= "0010101011100";
Trees_din <= "00000000010000010001011011001001";
wait for Clk_period;
Addr <= "0010101011101";
Trees_din <= "00000000000000000010010100001000";
wait for Clk_period;
Addr <= "0010101011110";
Trees_din <= "00000101000000000100011000000100";
wait for Clk_period;
Addr <= "0010101011111";
Trees_din <= "00000000001000100001011011001001";
wait for Clk_period;
Addr <= "0010101100000";
Trees_din <= "00000000010000000001011011001001";
wait for Clk_period;
Addr <= "0010101100001";
Trees_din <= "00000010000000000010010100000100";
wait for Clk_period;
Addr <= "0010101100010";
Trees_din <= "00000000010101100001011011001001";
wait for Clk_period;
Addr <= "0010101100011";
Trees_din <= "00000000000010010001011011001001";
wait for Clk_period;
Addr <= "0010101100100";
Trees_din <= "00000001000000000001001000010000";
wait for Clk_period;
Addr <= "0010101100101";
Trees_din <= "00000100000000000001111000001000";
wait for Clk_period;
Addr <= "0010101100110";
Trees_din <= "00000001000000000010010000000100";
wait for Clk_period;
Addr <= "0010101100111";
Trees_din <= "00000000010010110001011011001001";
wait for Clk_period;
Addr <= "0010101101000";
Trees_din <= "00000000010001000001011011001001";
wait for Clk_period;
Addr <= "0010101101001";
Trees_din <= "00000100000000000000101100000100";
wait for Clk_period;
Addr <= "0010101101010";
Trees_din <= "00000000010111000001011011001001";
wait for Clk_period;
Addr <= "0010101101011";
Trees_din <= "00000000001010000001011011001001";
wait for Clk_period;
Addr <= "0010101101100";
Trees_din <= "00000001000000000000001000001000";
wait for Clk_period;
Addr <= "0010101101101";
Trees_din <= "00000110000000000101100000000100";
wait for Clk_period;
Addr <= "0010101101110";
Trees_din <= "00000000001110110001011011001001";
wait for Clk_period;
Addr <= "0010101101111";
Trees_din <= "00000000001100110001011011001001";
wait for Clk_period;
Addr <= "0010101110000";
Trees_din <= "00000000000000000001100000000100";
wait for Clk_period;
Addr <= "0010101110001";
Trees_din <= "00000000001100100001011011001001";
wait for Clk_period;
Addr <= "0010101110010";
Trees_din <= "00000000000011110001011011001001";
wait for Clk_period;
Addr <= "0010101110011";
Trees_din <= "00000010000000000011101001000000";
wait for Clk_period;
Addr <= "0010101110100";
Trees_din <= "00000000000000000010110000100000";
wait for Clk_period;
Addr <= "0010101110101";
Trees_din <= "00000010000000000100000000010000";
wait for Clk_period;
Addr <= "0010101110110";
Trees_din <= "00000110000000000010010000001000";
wait for Clk_period;
Addr <= "0010101110111";
Trees_din <= "00000110000000000001001100000100";
wait for Clk_period;
Addr <= "0010101111000";
Trees_din <= "00000000000000110001011011001001";
wait for Clk_period;
Addr <= "0010101111001";
Trees_din <= "00000000000111000001011011001001";
wait for Clk_period;
Addr <= "0010101111010";
Trees_din <= "00000111000000000010001100000100";
wait for Clk_period;
Addr <= "0010101111011";
Trees_din <= "00000000000101100001011011001001";
wait for Clk_period;
Addr <= "0010101111100";
Trees_din <= "00000000010101100001011011001001";
wait for Clk_period;
Addr <= "0010101111101";
Trees_din <= "00000111000000000100001000001000";
wait for Clk_period;
Addr <= "0010101111110";
Trees_din <= "00000010000000000011111100000100";
wait for Clk_period;
Addr <= "0010101111111";
Trees_din <= "00000000001000100001011011001001";
wait for Clk_period;
Addr <= "0010110000000";
Trees_din <= "00000000000101100001011011001001";
wait for Clk_period;
Addr <= "0010110000001";
Trees_din <= "00000011000000000011100100000100";
wait for Clk_period;
Addr <= "0010110000010";
Trees_din <= "00000000011000100001011011001001";
wait for Clk_period;
Addr <= "0010110000011";
Trees_din <= "00000000000100010001011011001001";
wait for Clk_period;
Addr <= "0010110000100";
Trees_din <= "00000001000000000110001100010000";
wait for Clk_period;
Addr <= "0010110000101";
Trees_din <= "00000101000000000101011000001000";
wait for Clk_period;
Addr <= "0010110000110";
Trees_din <= "00000111000000000101111100000100";
wait for Clk_period;
Addr <= "0010110000111";
Trees_din <= "00000000010101000001011011001001";
wait for Clk_period;
Addr <= "0010110001000";
Trees_din <= "00000000010111000001011011001001";
wait for Clk_period;
Addr <= "0010110001001";
Trees_din <= "00000010000000000110001100000100";
wait for Clk_period;
Addr <= "0010110001010";
Trees_din <= "00000000000110010001011011001001";
wait for Clk_period;
Addr <= "0010110001011";
Trees_din <= "00000000010000000001011011001001";
wait for Clk_period;
Addr <= "0010110001100";
Trees_din <= "00000000000000000010100000001000";
wait for Clk_period;
Addr <= "0010110001101";
Trees_din <= "00000100000000000011000100000100";
wait for Clk_period;
Addr <= "0010110001110";
Trees_din <= "00000000001111100001011011001001";
wait for Clk_period;
Addr <= "0010110001111";
Trees_din <= "00000000001111000001011011001001";
wait for Clk_period;
Addr <= "0010110010000";
Trees_din <= "00000100000000000010010000000100";
wait for Clk_period;
Addr <= "0010110010001";
Trees_din <= "00000000010000000001011011001001";
wait for Clk_period;
Addr <= "0010110010010";
Trees_din <= "00000000010100010001011011001001";
wait for Clk_period;
Addr <= "0010110010011";
Trees_din <= "00000110000000000100100000100000";
wait for Clk_period;
Addr <= "0010110010100";
Trees_din <= "00000000000000000101011000010000";
wait for Clk_period;
Addr <= "0010110010101";
Trees_din <= "00000010000000000011001100001000";
wait for Clk_period;
Addr <= "0010110010110";
Trees_din <= "00000000000000000001111000000100";
wait for Clk_period;
Addr <= "0010110010111";
Trees_din <= "00000000001010000001011011001001";
wait for Clk_period;
Addr <= "0010110011000";
Trees_din <= "00000000011000000001011011001001";
wait for Clk_period;
Addr <= "0010110011001";
Trees_din <= "00000011000000000010100100000100";
wait for Clk_period;
Addr <= "0010110011010";
Trees_din <= "00000000010011110001011011001001";
wait for Clk_period;
Addr <= "0010110011011";
Trees_din <= "00000000000010110001011011001001";
wait for Clk_period;
Addr <= "0010110011100";
Trees_din <= "00000101000000000001000000001000";
wait for Clk_period;
Addr <= "0010110011101";
Trees_din <= "00000000000000000011110000000100";
wait for Clk_period;
Addr <= "0010110011110";
Trees_din <= "00000000000000110001011011001001";
wait for Clk_period;
Addr <= "0010110011111";
Trees_din <= "00000000001001100001011011001001";
wait for Clk_period;
Addr <= "0010110100000";
Trees_din <= "00000101000000000000101100000100";
wait for Clk_period;
Addr <= "0010110100001";
Trees_din <= "00000000000010000001011011001001";
wait for Clk_period;
Addr <= "0010110100010";
Trees_din <= "00000000001110000001011011001001";
wait for Clk_period;
Addr <= "0010110100011";
Trees_din <= "00000000000000000010010000010000";
wait for Clk_period;
Addr <= "0010110100100";
Trees_din <= "00000101000000000001111100001000";
wait for Clk_period;
Addr <= "0010110100101";
Trees_din <= "00000110000000000100101100000100";
wait for Clk_period;
Addr <= "0010110100110";
Trees_din <= "00000000010001110001011011001001";
wait for Clk_period;
Addr <= "0010110100111";
Trees_din <= "00000000000001100001011011001001";
wait for Clk_period;
Addr <= "0010110101000";
Trees_din <= "00000000000000000001011000000100";
wait for Clk_period;
Addr <= "0010110101001";
Trees_din <= "00000000001000100001011011001001";
wait for Clk_period;
Addr <= "0010110101010";
Trees_din <= "00000000000101110001011011001001";
wait for Clk_period;
Addr <= "0010110101011";
Trees_din <= "00000001000000000010100000001000";
wait for Clk_period;
Addr <= "0010110101100";
Trees_din <= "00000101000000000011010100000100";
wait for Clk_period;
Addr <= "0010110101101";
Trees_din <= "00000000001001010001011011001001";
wait for Clk_period;
Addr <= "0010110101110";
Trees_din <= "00000000001111010001011011001001";
wait for Clk_period;
Addr <= "0010110101111";
Trees_din <= "00000011000000000001011000000100";
wait for Clk_period;
Addr <= "0010110110000";
Trees_din <= "00000000000010000001011011001001";
wait for Clk_period;
Addr <= "0010110110001";
Trees_din <= "00000000001111010001011011001001";
wait for Clk_period;



----------tree 11-------------------

Addr <= "0010110110010";
Trees_din <= "00000010000000000000111010000000";
wait for Clk_period;
Addr <= "0010110110011";
Trees_din <= "00000111000000000101101001000000";
wait for Clk_period;
Addr <= "0010110110100";
Trees_din <= "00000111000000000010110100100000";
wait for Clk_period;
Addr <= "0010110110101";
Trees_din <= "00000110000000000011000100010000";
wait for Clk_period;
Addr <= "0010110110110";
Trees_din <= "00000001000000000001010000001000";
wait for Clk_period;
Addr <= "0010110110111";
Trees_din <= "00000101000000000100110100000100";
wait for Clk_period;
Addr <= "0010110111000";
Trees_din <= "00000000010001010001100011000101";
wait for Clk_period;
Addr <= "0010110111001";
Trees_din <= "00000000001010110001100011000101";
wait for Clk_period;
Addr <= "0010110111010";
Trees_din <= "00000111000000000011000000000100";
wait for Clk_period;
Addr <= "0010110111011";
Trees_din <= "00000000000111110001100011000101";
wait for Clk_period;
Addr <= "0010110111100";
Trees_din <= "00000000001001100001100011000101";
wait for Clk_period;
Addr <= "0010110111101";
Trees_din <= "00000100000000000110000000001000";
wait for Clk_period;
Addr <= "0010110111110";
Trees_din <= "00000110000000000110001000000100";
wait for Clk_period;
Addr <= "0010110111111";
Trees_din <= "00000000011000010001100011000101";
wait for Clk_period;
Addr <= "0010111000000";
Trees_din <= "00000000001100110001100011000101";
wait for Clk_period;
Addr <= "0010111000001";
Trees_din <= "00000111000000000011011000000100";
wait for Clk_period;
Addr <= "0010111000010";
Trees_din <= "00000000000100100001100011000101";
wait for Clk_period;
Addr <= "0010111000011";
Trees_din <= "00000000010010000001100011000101";
wait for Clk_period;
Addr <= "0010111000100";
Trees_din <= "00000011000000000000100000010000";
wait for Clk_period;
Addr <= "0010111000101";
Trees_din <= "00000100000000000110001000001000";
wait for Clk_period;
Addr <= "0010111000110";
Trees_din <= "00000111000000000010101000000100";
wait for Clk_period;
Addr <= "0010111000111";
Trees_din <= "00000000000111100001100011000101";
wait for Clk_period;
Addr <= "0010111001000";
Trees_din <= "00000000010100000001100011000101";
wait for Clk_period;
Addr <= "0010111001001";
Trees_din <= "00000011000000000100100000000100";
wait for Clk_period;
Addr <= "0010111001010";
Trees_din <= "00000000000010100001100011000101";
wait for Clk_period;
Addr <= "0010111001011";
Trees_din <= "00000000000100000001100011000101";
wait for Clk_period;
Addr <= "0010111001100";
Trees_din <= "00000101000000000101001100001000";
wait for Clk_period;
Addr <= "0010111001101";
Trees_din <= "00000011000000000100110100000100";
wait for Clk_period;
Addr <= "0010111001110";
Trees_din <= "00000000001001000001100011000101";
wait for Clk_period;
Addr <= "0010111001111";
Trees_din <= "00000000010000000001100011000101";
wait for Clk_period;
Addr <= "0010111010000";
Trees_din <= "00000110000000000001001100000100";
wait for Clk_period;
Addr <= "0010111010001";
Trees_din <= "00000000010011100001100011000101";
wait for Clk_period;
Addr <= "0010111010010";
Trees_din <= "00000000001100010001100011000101";
wait for Clk_period;
Addr <= "0010111010011";
Trees_din <= "00000110000000000001011000100000";
wait for Clk_period;
Addr <= "0010111010100";
Trees_din <= "00000001000000000100000000010000";
wait for Clk_period;
Addr <= "0010111010101";
Trees_din <= "00000010000000000101100100001000";
wait for Clk_period;
Addr <= "0010111010110";
Trees_din <= "00000110000000000010000000000100";
wait for Clk_period;
Addr <= "0010111010111";
Trees_din <= "00000000001111010001100011000101";
wait for Clk_period;
Addr <= "0010111011000";
Trees_din <= "00000000001101000001100011000101";
wait for Clk_period;
Addr <= "0010111011001";
Trees_din <= "00000101000000000011011100000100";
wait for Clk_period;
Addr <= "0010111011010";
Trees_din <= "00000000010000110001100011000101";
wait for Clk_period;
Addr <= "0010111011011";
Trees_din <= "00000000000111000001100011000101";
wait for Clk_period;
Addr <= "0010111011100";
Trees_din <= "00000001000000000101110000001000";
wait for Clk_period;
Addr <= "0010111011101";
Trees_din <= "00000010000000000011001100000100";
wait for Clk_period;
Addr <= "0010111011110";
Trees_din <= "00000000010100110001100011000101";
wait for Clk_period;
Addr <= "0010111011111";
Trees_din <= "00000000000011000001100011000101";
wait for Clk_period;
Addr <= "0010111100000";
Trees_din <= "00000001000000000001010100000100";
wait for Clk_period;
Addr <= "0010111100001";
Trees_din <= "00000000001111000001100011000101";
wait for Clk_period;
Addr <= "0010111100010";
Trees_din <= "00000000001001100001100011000101";
wait for Clk_period;
Addr <= "0010111100011";
Trees_din <= "00000111000000000011100000010000";
wait for Clk_period;
Addr <= "0010111100100";
Trees_din <= "00000010000000000001010100001000";
wait for Clk_period;
Addr <= "0010111100101";
Trees_din <= "00000010000000000011010000000100";
wait for Clk_period;
Addr <= "0010111100110";
Trees_din <= "00000000011000010001100011000101";
wait for Clk_period;
Addr <= "0010111100111";
Trees_din <= "00000000010011010001100011000101";
wait for Clk_period;
Addr <= "0010111101000";
Trees_din <= "00000001000000000000001000000100";
wait for Clk_period;
Addr <= "0010111101001";
Trees_din <= "00000000000001100001100011000101";
wait for Clk_period;
Addr <= "0010111101010";
Trees_din <= "00000000001000110001100011000101";
wait for Clk_period;
Addr <= "0010111101011";
Trees_din <= "00000100000000000100001100001000";
wait for Clk_period;
Addr <= "0010111101100";
Trees_din <= "00000100000000000100101000000100";
wait for Clk_period;
Addr <= "0010111101101";
Trees_din <= "00000000000000000001100011000101";
wait for Clk_period;
Addr <= "0010111101110";
Trees_din <= "00000000000000000001100011000101";
wait for Clk_period;
Addr <= "0010111101111";
Trees_din <= "00000110000000000001011100000100";
wait for Clk_period;
Addr <= "0010111110000";
Trees_din <= "00000000010001000001100011000101";
wait for Clk_period;
Addr <= "0010111110001";
Trees_din <= "00000000000110110001100011000101";
wait for Clk_period;
Addr <= "0010111110010";
Trees_din <= "00000111000000000010010101000000";
wait for Clk_period;
Addr <= "0010111110011";
Trees_din <= "00000100000000000011100000100000";
wait for Clk_period;
Addr <= "0010111110100";
Trees_din <= "00000100000000000100111100010000";
wait for Clk_period;
Addr <= "0010111110101";
Trees_din <= "00000101000000000001101000001000";
wait for Clk_period;
Addr <= "0010111110110";
Trees_din <= "00000000000000000011100000000100";
wait for Clk_period;
Addr <= "0010111110111";
Trees_din <= "00000000010001010001100011000101";
wait for Clk_period;
Addr <= "0010111111000";
Trees_din <= "00000000000101010001100011000101";
wait for Clk_period;
Addr <= "0010111111001";
Trees_din <= "00000001000000000010000100000100";
wait for Clk_period;
Addr <= "0010111111010";
Trees_din <= "00000000010111010001100011000101";
wait for Clk_period;
Addr <= "0010111111011";
Trees_din <= "00000000001100010001100011000101";
wait for Clk_period;
Addr <= "0010111111100";
Trees_din <= "00000010000000000100110100001000";
wait for Clk_period;
Addr <= "0010111111101";
Trees_din <= "00000101000000000101001000000100";
wait for Clk_period;
Addr <= "0010111111110";
Trees_din <= "00000000010101000001100011000101";
wait for Clk_period;
Addr <= "0010111111111";
Trees_din <= "00000000000000110001100011000101";
wait for Clk_period;
Addr <= "0011000000000";
Trees_din <= "00000111000000000010110100000100";
wait for Clk_period;
Addr <= "0011000000001";
Trees_din <= "00000000000010100001100011000101";
wait for Clk_period;
Addr <= "0011000000010";
Trees_din <= "00000000001101000001100011000101";
wait for Clk_period;
Addr <= "0011000000011";
Trees_din <= "00000001000000000100011000010000";
wait for Clk_period;
Addr <= "0011000000100";
Trees_din <= "00000100000000000100100100001000";
wait for Clk_period;
Addr <= "0011000000101";
Trees_din <= "00000110000000000100101100000100";
wait for Clk_period;
Addr <= "0011000000110";
Trees_din <= "00000000010101100001100011000101";
wait for Clk_period;
Addr <= "0011000000111";
Trees_din <= "00000000001011000001100011000101";
wait for Clk_period;
Addr <= "0011000001000";
Trees_din <= "00000000000000000011000000000100";
wait for Clk_period;
Addr <= "0011000001001";
Trees_din <= "00000000010011110001100011000101";
wait for Clk_period;
Addr <= "0011000001010";
Trees_din <= "00000000000100100001100011000101";
wait for Clk_period;
Addr <= "0011000001011";
Trees_din <= "00000111000000000001000100001000";
wait for Clk_period;
Addr <= "0011000001100";
Trees_din <= "00000111000000000101011000000100";
wait for Clk_period;
Addr <= "0011000001101";
Trees_din <= "00000000001010110001100011000101";
wait for Clk_period;
Addr <= "0011000001110";
Trees_din <= "00000000001000010001100011000101";
wait for Clk_period;
Addr <= "0011000001111";
Trees_din <= "00000001000000000101111000000100";
wait for Clk_period;
Addr <= "0011000010000";
Trees_din <= "00000000000001110001100011000101";
wait for Clk_period;
Addr <= "0011000010001";
Trees_din <= "00000000010111110001100011000101";
wait for Clk_period;
Addr <= "0011000010010";
Trees_din <= "00000111000000000100101000100000";
wait for Clk_period;
Addr <= "0011000010011";
Trees_din <= "00000100000000000101010100010000";
wait for Clk_period;
Addr <= "0011000010100";
Trees_din <= "00000001000000000001011100001000";
wait for Clk_period;
Addr <= "0011000010101";
Trees_din <= "00000011000000000110000000000100";
wait for Clk_period;
Addr <= "0011000010110";
Trees_din <= "00000000010011100001100011000101";
wait for Clk_period;
Addr <= "0011000010111";
Trees_din <= "00000000001011100001100011000101";
wait for Clk_period;
Addr <= "0011000011000";
Trees_din <= "00000101000000000100111100000100";
wait for Clk_period;
Addr <= "0011000011001";
Trees_din <= "00000000000011110001100011000101";
wait for Clk_period;
Addr <= "0011000011010";
Trees_din <= "00000000001010000001100011000101";
wait for Clk_period;
Addr <= "0011000011011";
Trees_din <= "00000001000000000010001000001000";
wait for Clk_period;
Addr <= "0011000011100";
Trees_din <= "00000110000000000011100100000100";
wait for Clk_period;
Addr <= "0011000011101";
Trees_din <= "00000000010100000001100011000101";
wait for Clk_period;
Addr <= "0011000011110";
Trees_din <= "00000000001110010001100011000101";
wait for Clk_period;
Addr <= "0011000011111";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "0011000100000";
Trees_din <= "00000000001111100001100011000101";
wait for Clk_period;
Addr <= "0011000100001";
Trees_din <= "00000000000101000001100011000101";
wait for Clk_period;
Addr <= "0011000100010";
Trees_din <= "00000000000000000010000100010000";
wait for Clk_period;
Addr <= "0011000100011";
Trees_din <= "00000001000000000101010000001000";
wait for Clk_period;
Addr <= "0011000100100";
Trees_din <= "00000011000000000110000100000100";
wait for Clk_period;
Addr <= "0011000100101";
Trees_din <= "00000000001001100001100011000101";
wait for Clk_period;
Addr <= "0011000100110";
Trees_din <= "00000000010000010001100011000101";
wait for Clk_period;
Addr <= "0011000100111";
Trees_din <= "00000100000000000011110100000100";
wait for Clk_period;
Addr <= "0011000101000";
Trees_din <= "00000000010110110001100011000101";
wait for Clk_period;
Addr <= "0011000101001";
Trees_din <= "00000000010111100001100011000101";
wait for Clk_period;
Addr <= "0011000101010";
Trees_din <= "00000111000000000010011100001000";
wait for Clk_period;
Addr <= "0011000101011";
Trees_din <= "00000011000000000001001100000100";
wait for Clk_period;
Addr <= "0011000101100";
Trees_din <= "00000000000110100001100011000101";
wait for Clk_period;
Addr <= "0011000101101";
Trees_din <= "00000000010010000001100011000101";
wait for Clk_period;
Addr <= "0011000101110";
Trees_din <= "00000110000000000011010100000100";
wait for Clk_period;
Addr <= "0011000101111";
Trees_din <= "00000000001000000001100011000101";
wait for Clk_period;
Addr <= "0011000110000";
Trees_din <= "00000000010010000001100011000101";
wait for Clk_period;



----------tree 12-------------------

Addr <= "0011000110001";
Trees_din <= "00000011000000000011011110000000";
wait for Clk_period;
Addr <= "0011000110010";
Trees_din <= "00000111000000000101001001000000";
wait for Clk_period;
Addr <= "0011000110011";
Trees_din <= "00000011000000000100011100100000";
wait for Clk_period;
Addr <= "0011000110100";
Trees_din <= "00000011000000000000100100010000";
wait for Clk_period;
Addr <= "0011000110101";
Trees_din <= "00000111000000000010100100001000";
wait for Clk_period;
Addr <= "0011000110110";
Trees_din <= "00000010000000000010111000000100";
wait for Clk_period;
Addr <= "0011000110111";
Trees_din <= "00000000000101110001101011000001";
wait for Clk_period;
Addr <= "0011000111000";
Trees_din <= "00000000001111110001101011000001";
wait for Clk_period;
Addr <= "0011000111001";
Trees_din <= "00000110000000000011010100000100";
wait for Clk_period;
Addr <= "0011000111010";
Trees_din <= "00000000010100010001101011000001";
wait for Clk_period;
Addr <= "0011000111011";
Trees_din <= "00000000001011110001101011000001";
wait for Clk_period;
Addr <= "0011000111100";
Trees_din <= "00000010000000000011000100001000";
wait for Clk_period;
Addr <= "0011000111101";
Trees_din <= "00000001000000000000111000000100";
wait for Clk_period;
Addr <= "0011000111110";
Trees_din <= "00000000010111110001101011000001";
wait for Clk_period;
Addr <= "0011000111111";
Trees_din <= "00000000001011100001101011000001";
wait for Clk_period;
Addr <= "0011001000000";
Trees_din <= "00000010000000000010111000000100";
wait for Clk_period;
Addr <= "0011001000001";
Trees_din <= "00000000001010000001101011000001";
wait for Clk_period;
Addr <= "0011001000010";
Trees_din <= "00000000000111010001101011000001";
wait for Clk_period;
Addr <= "0011001000011";
Trees_din <= "00000101000000000010111100010000";
wait for Clk_period;
Addr <= "0011001000100";
Trees_din <= "00000100000000000100000100001000";
wait for Clk_period;
Addr <= "0011001000101";
Trees_din <= "00000101000000000100011100000100";
wait for Clk_period;
Addr <= "0011001000110";
Trees_din <= "00000000001000100001101011000001";
wait for Clk_period;
Addr <= "0011001000111";
Trees_din <= "00000000001000110001101011000001";
wait for Clk_period;
Addr <= "0011001001000";
Trees_din <= "00000100000000000001011000000100";
wait for Clk_period;
Addr <= "0011001001001";
Trees_din <= "00000000010011110001101011000001";
wait for Clk_period;
Addr <= "0011001001010";
Trees_din <= "00000000010001110001101011000001";
wait for Clk_period;
Addr <= "0011001001011";
Trees_din <= "00000101000000000000110000001000";
wait for Clk_period;
Addr <= "0011001001100";
Trees_din <= "00000101000000000011001000000100";
wait for Clk_period;
Addr <= "0011001001101";
Trees_din <= "00000000010110000001101011000001";
wait for Clk_period;
Addr <= "0011001001110";
Trees_din <= "00000000010111100001101011000001";
wait for Clk_period;
Addr <= "0011001001111";
Trees_din <= "00000011000000000001011100000100";
wait for Clk_period;
Addr <= "0011001010000";
Trees_din <= "00000000000010110001101011000001";
wait for Clk_period;
Addr <= "0011001010001";
Trees_din <= "00000000010011010001101011000001";
wait for Clk_period;
Addr <= "0011001010010";
Trees_din <= "00000111000000000000010000100000";
wait for Clk_period;
Addr <= "0011001010011";
Trees_din <= "00000011000000000011000100010000";
wait for Clk_period;
Addr <= "0011001010100";
Trees_din <= "00000100000000000100110100001000";
wait for Clk_period;
Addr <= "0011001010101";
Trees_din <= "00000101000000000011011100000100";
wait for Clk_period;
Addr <= "0011001010110";
Trees_din <= "00000000010011010001101011000001";
wait for Clk_period;
Addr <= "0011001010111";
Trees_din <= "00000000010100000001101011000001";
wait for Clk_period;
Addr <= "0011001011000";
Trees_din <= "00000001000000000101010000000100";
wait for Clk_period;
Addr <= "0011001011001";
Trees_din <= "00000000010010100001101011000001";
wait for Clk_period;
Addr <= "0011001011010";
Trees_din <= "00000000000111100001101011000001";
wait for Clk_period;
Addr <= "0011001011011";
Trees_din <= "00000110000000000101111100001000";
wait for Clk_period;
Addr <= "0011001011100";
Trees_din <= "00000011000000000100101100000100";
wait for Clk_period;
Addr <= "0011001011101";
Trees_din <= "00000000010011000001101011000001";
wait for Clk_period;
Addr <= "0011001011110";
Trees_din <= "00000000000100100001101011000001";
wait for Clk_period;
Addr <= "0011001011111";
Trees_din <= "00000110000000000000110100000100";
wait for Clk_period;
Addr <= "0011001100000";
Trees_din <= "00000000010010100001101011000001";
wait for Clk_period;
Addr <= "0011001100001";
Trees_din <= "00000000001000100001101011000001";
wait for Clk_period;
Addr <= "0011001100010";
Trees_din <= "00000111000000000010110000010000";
wait for Clk_period;
Addr <= "0011001100011";
Trees_din <= "00000001000000000110000100001000";
wait for Clk_period;
Addr <= "0011001100100";
Trees_din <= "00000010000000000001100100000100";
wait for Clk_period;
Addr <= "0011001100101";
Trees_din <= "00000000001000110001101011000001";
wait for Clk_period;
Addr <= "0011001100110";
Trees_din <= "00000000010100110001101011000001";
wait for Clk_period;
Addr <= "0011001100111";
Trees_din <= "00000010000000000001110000000100";
wait for Clk_period;
Addr <= "0011001101000";
Trees_din <= "00000000000000000001101011000001";
wait for Clk_period;
Addr <= "0011001101001";
Trees_din <= "00000000001011110001101011000001";
wait for Clk_period;
Addr <= "0011001101010";
Trees_din <= "00000011000000000100100000001000";
wait for Clk_period;
Addr <= "0011001101011";
Trees_din <= "00000010000000000010100100000100";
wait for Clk_period;
Addr <= "0011001101100";
Trees_din <= "00000000000010110001101011000001";
wait for Clk_period;
Addr <= "0011001101101";
Trees_din <= "00000000000001100001101011000001";
wait for Clk_period;
Addr <= "0011001101110";
Trees_din <= "00000111000000000101011100000100";
wait for Clk_period;
Addr <= "0011001101111";
Trees_din <= "00000000010011010001101011000001";
wait for Clk_period;
Addr <= "0011001110000";
Trees_din <= "00000000000000110001101011000001";
wait for Clk_period;
Addr <= "0011001110001";
Trees_din <= "00000010000000000001100101000000";
wait for Clk_period;
Addr <= "0011001110010";
Trees_din <= "00000110000000000011011000100000";
wait for Clk_period;
Addr <= "0011001110011";
Trees_din <= "00000010000000000011000000010000";
wait for Clk_period;
Addr <= "0011001110100";
Trees_din <= "00000110000000000100111000001000";
wait for Clk_period;
Addr <= "0011001110101";
Trees_din <= "00000111000000000010010100000100";
wait for Clk_period;
Addr <= "0011001110110";
Trees_din <= "00000000010100000001101011000001";
wait for Clk_period;
Addr <= "0011001110111";
Trees_din <= "00000000000001100001101011000001";
wait for Clk_period;
Addr <= "0011001111000";
Trees_din <= "00000101000000000011100100000100";
wait for Clk_period;
Addr <= "0011001111001";
Trees_din <= "00000000010111100001101011000001";
wait for Clk_period;
Addr <= "0011001111010";
Trees_din <= "00000000010011100001101011000001";
wait for Clk_period;
Addr <= "0011001111011";
Trees_din <= "00000001000000000000010000001000";
wait for Clk_period;
Addr <= "0011001111100";
Trees_din <= "00000011000000000000000000000100";
wait for Clk_period;
Addr <= "0011001111101";
Trees_din <= "00000000001111000001101011000001";
wait for Clk_period;
Addr <= "0011001111110";
Trees_din <= "00000000001001010001101011000001";
wait for Clk_period;
Addr <= "0011001111111";
Trees_din <= "00000100000000000100001000000100";
wait for Clk_period;
Addr <= "0011010000000";
Trees_din <= "00000000000001000001101011000001";
wait for Clk_period;
Addr <= "0011010000001";
Trees_din <= "00000000010111000001101011000001";
wait for Clk_period;
Addr <= "0011010000010";
Trees_din <= "00000001000000000010011000010000";
wait for Clk_period;
Addr <= "0011010000011";
Trees_din <= "00000000000000000011110000001000";
wait for Clk_period;
Addr <= "0011010000100";
Trees_din <= "00000110000000000100111100000100";
wait for Clk_period;
Addr <= "0011010000101";
Trees_din <= "00000000000011000001101011000001";
wait for Clk_period;
Addr <= "0011010000110";
Trees_din <= "00000000001101100001101011000001";
wait for Clk_period;
Addr <= "0011010000111";
Trees_din <= "00000000000000000100001000000100";
wait for Clk_period;
Addr <= "0011010001000";
Trees_din <= "00000000001101110001101011000001";
wait for Clk_period;
Addr <= "0011010001001";
Trees_din <= "00000000000011000001101011000001";
wait for Clk_period;
Addr <= "0011010001010";
Trees_din <= "00000011000000000001001000001000";
wait for Clk_period;
Addr <= "0011010001011";
Trees_din <= "00000000000000000011010100000100";
wait for Clk_period;
Addr <= "0011010001100";
Trees_din <= "00000000001001010001101011000001";
wait for Clk_period;
Addr <= "0011010001101";
Trees_din <= "00000000010100110001101011000001";
wait for Clk_period;
Addr <= "0011010001110";
Trees_din <= "00000111000000000101011100000100";
wait for Clk_period;
Addr <= "0011010001111";
Trees_din <= "00000000010111000001101011000001";
wait for Clk_period;
Addr <= "0011010010000";
Trees_din <= "00000000000011000001101011000001";
wait for Clk_period;
Addr <= "0011010010001";
Trees_din <= "00000000000000000010111100100000";
wait for Clk_period;
Addr <= "0011010010010";
Trees_din <= "00000011000000000011101000010000";
wait for Clk_period;
Addr <= "0011010010011";
Trees_din <= "00000001000000000101101100001000";
wait for Clk_period;
Addr <= "0011010010100";
Trees_din <= "00000101000000000010110100000100";
wait for Clk_period;
Addr <= "0011010010101";
Trees_din <= "00000000000011000001101011000001";
wait for Clk_period;
Addr <= "0011010010110";
Trees_din <= "00000000000010000001101011000001";
wait for Clk_period;
Addr <= "0011010010111";
Trees_din <= "00000000000000000010001000000100";
wait for Clk_period;
Addr <= "0011010011000";
Trees_din <= "00000000010000110001101011000001";
wait for Clk_period;
Addr <= "0011010011001";
Trees_din <= "00000000010010100001101011000001";
wait for Clk_period;
Addr <= "0011010011010";
Trees_din <= "00000011000000000001100100001000";
wait for Clk_period;
Addr <= "0011010011011";
Trees_din <= "00000010000000000011110100000100";
wait for Clk_period;
Addr <= "0011010011100";
Trees_din <= "00000000000011100001101011000001";
wait for Clk_period;
Addr <= "0011010011101";
Trees_din <= "00000000000101100001101011000001";
wait for Clk_period;
Addr <= "0011010011110";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "0011010011111";
Trees_din <= "00000000001110010001101011000001";
wait for Clk_period;
Addr <= "0011010100000";
Trees_din <= "00000000000110000001101011000001";
wait for Clk_period;
Addr <= "0011010100001";
Trees_din <= "00000100000000000000010100010000";
wait for Clk_period;
Addr <= "0011010100010";
Trees_din <= "00000001000000000010110000001000";
wait for Clk_period;
Addr <= "0011010100011";
Trees_din <= "00000011000000000100000100000100";
wait for Clk_period;
Addr <= "0011010100100";
Trees_din <= "00000000010100110001101011000001";
wait for Clk_period;
Addr <= "0011010100101";
Trees_din <= "00000000000011010001101011000001";
wait for Clk_period;
Addr <= "0011010100110";
Trees_din <= "00000110000000000010001100000100";
wait for Clk_period;
Addr <= "0011010100111";
Trees_din <= "00000000001011010001101011000001";
wait for Clk_period;
Addr <= "0011010101000";
Trees_din <= "00000000000111110001101011000001";
wait for Clk_period;
Addr <= "0011010101001";
Trees_din <= "00000110000000000100101100001000";
wait for Clk_period;
Addr <= "0011010101010";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "0011010101011";
Trees_din <= "00000000010001110001101011000001";
wait for Clk_period;
Addr <= "0011010101100";
Trees_din <= "00000000001110000001101011000001";
wait for Clk_period;
Addr <= "0011010101101";
Trees_din <= "00000110000000000010000000000100";
wait for Clk_period;
Addr <= "0011010101110";
Trees_din <= "00000000001000100001101011000001";
wait for Clk_period;
Addr <= "0011010101111";
Trees_din <= "00000000000101010001101011000001";
wait for Clk_period;



----------tree 13-------------------

Addr <= "0011010110000";
Trees_din <= "00000110000000000100101010000000";
wait for Clk_period;
Addr <= "0011010110001";
Trees_din <= "00000010000000000100100101000000";
wait for Clk_period;
Addr <= "0011010110010";
Trees_din <= "00000101000000000101111100100000";
wait for Clk_period;
Addr <= "0011010110011";
Trees_din <= "00000011000000000011010000010000";
wait for Clk_period;
Addr <= "0011010110100";
Trees_din <= "00000010000000000001010000001000";
wait for Clk_period;
Addr <= "0011010110101";
Trees_din <= "00000111000000000001111100000100";
wait for Clk_period;
Addr <= "0011010110110";
Trees_din <= "00000000000010110001110010111101";
wait for Clk_period;
Addr <= "0011010110111";
Trees_din <= "00000000001110100001110010111101";
wait for Clk_period;
Addr <= "0011010111000";
Trees_din <= "00000011000000000010011100000100";
wait for Clk_period;
Addr <= "0011010111001";
Trees_din <= "00000000000000100001110010111101";
wait for Clk_period;
Addr <= "0011010111010";
Trees_din <= "00000000001101000001110010111101";
wait for Clk_period;
Addr <= "0011010111011";
Trees_din <= "00000101000000000001001000001000";
wait for Clk_period;
Addr <= "0011010111100";
Trees_din <= "00000101000000000011100000000100";
wait for Clk_period;
Addr <= "0011010111101";
Trees_din <= "00000000010101110001110010111101";
wait for Clk_period;
Addr <= "0011010111110";
Trees_din <= "00000000010110110001110010111101";
wait for Clk_period;
Addr <= "0011010111111";
Trees_din <= "00000001000000000000010000000100";
wait for Clk_period;
Addr <= "0011011000000";
Trees_din <= "00000000001110110001110010111101";
wait for Clk_period;
Addr <= "0011011000001";
Trees_din <= "00000000001100100001110010111101";
wait for Clk_period;
Addr <= "0011011000010";
Trees_din <= "00000000000000000101010100010000";
wait for Clk_period;
Addr <= "0011011000011";
Trees_din <= "00000101000000000010101000001000";
wait for Clk_period;
Addr <= "0011011000100";
Trees_din <= "00000110000000000000010100000100";
wait for Clk_period;
Addr <= "0011011000101";
Trees_din <= "00000000001101100001110010111101";
wait for Clk_period;
Addr <= "0011011000110";
Trees_din <= "00000000010010100001110010111101";
wait for Clk_period;
Addr <= "0011011000111";
Trees_din <= "00000111000000000000011100000100";
wait for Clk_period;
Addr <= "0011011001000";
Trees_din <= "00000000011001000001110010111101";
wait for Clk_period;
Addr <= "0011011001001";
Trees_din <= "00000000001111100001110010111101";
wait for Clk_period;
Addr <= "0011011001010";
Trees_din <= "00000101000000000011000000001000";
wait for Clk_period;
Addr <= "0011011001011";
Trees_din <= "00000000000000000011000100000100";
wait for Clk_period;
Addr <= "0011011001100";
Trees_din <= "00000000001110000001110010111101";
wait for Clk_period;
Addr <= "0011011001101";
Trees_din <= "00000000001000110001110010111101";
wait for Clk_period;
Addr <= "0011011001110";
Trees_din <= "00000110000000000011010100000100";
wait for Clk_period;
Addr <= "0011011001111";
Trees_din <= "00000000001111000001110010111101";
wait for Clk_period;
Addr <= "0011011010000";
Trees_din <= "00000000000111100001110010111101";
wait for Clk_period;
Addr <= "0011011010001";
Trees_din <= "00000111000000000011000100100000";
wait for Clk_period;
Addr <= "0011011010010";
Trees_din <= "00000001000000000101000100010000";
wait for Clk_period;
Addr <= "0011011010011";
Trees_din <= "00000011000000000000110100001000";
wait for Clk_period;
Addr <= "0011011010100";
Trees_din <= "00000010000000000001001100000100";
wait for Clk_period;
Addr <= "0011011010101";
Trees_din <= "00000000000000000001110010111101";
wait for Clk_period;
Addr <= "0011011010110";
Trees_din <= "00000000000101010001110010111101";
wait for Clk_period;
Addr <= "0011011010111";
Trees_din <= "00000000000000000010010000000100";
wait for Clk_period;
Addr <= "0011011011000";
Trees_din <= "00000000010111110001110010111101";
wait for Clk_period;
Addr <= "0011011011001";
Trees_din <= "00000000011000110001110010111101";
wait for Clk_period;
Addr <= "0011011011010";
Trees_din <= "00000000000000000000010000001000";
wait for Clk_period;
Addr <= "0011011011011";
Trees_din <= "00000000000000000001101000000100";
wait for Clk_period;
Addr <= "0011011011100";
Trees_din <= "00000000000110110001110010111101";
wait for Clk_period;
Addr <= "0011011011101";
Trees_din <= "00000000000001000001110010111101";
wait for Clk_period;
Addr <= "0011011011110";
Trees_din <= "00000000000000000000011000000100";
wait for Clk_period;
Addr <= "0011011011111";
Trees_din <= "00000000000010000001110010111101";
wait for Clk_period;
Addr <= "0011011100000";
Trees_din <= "00000000010100000001110010111101";
wait for Clk_period;
Addr <= "0011011100001";
Trees_din <= "00000010000000000100100100010000";
wait for Clk_period;
Addr <= "0011011100010";
Trees_din <= "00000101000000000101101000001000";
wait for Clk_period;
Addr <= "0011011100011";
Trees_din <= "00000001000000000000100000000100";
wait for Clk_period;
Addr <= "0011011100100";
Trees_din <= "00000000010000010001110010111101";
wait for Clk_period;
Addr <= "0011011100101";
Trees_din <= "00000000001000100001110010111101";
wait for Clk_period;
Addr <= "0011011100110";
Trees_din <= "00000101000000000101100000000100";
wait for Clk_period;
Addr <= "0011011100111";
Trees_din <= "00000000000000010001110010111101";
wait for Clk_period;
Addr <= "0011011101000";
Trees_din <= "00000000010000010001110010111101";
wait for Clk_period;
Addr <= "0011011101001";
Trees_din <= "00000001000000000010001100001000";
wait for Clk_period;
Addr <= "0011011101010";
Trees_din <= "00000001000000000101100000000100";
wait for Clk_period;
Addr <= "0011011101011";
Trees_din <= "00000000010010100001110010111101";
wait for Clk_period;
Addr <= "0011011101100";
Trees_din <= "00000000010000110001110010111101";
wait for Clk_period;
Addr <= "0011011101101";
Trees_din <= "00000011000000000010001100000100";
wait for Clk_period;
Addr <= "0011011101110";
Trees_din <= "00000000000111000001110010111101";
wait for Clk_period;
Addr <= "0011011101111";
Trees_din <= "00000000001101010001110010111101";
wait for Clk_period;
Addr <= "0011011110000";
Trees_din <= "00000001000000000010011001000000";
wait for Clk_period;
Addr <= "0011011110001";
Trees_din <= "00000110000000000101000000100000";
wait for Clk_period;
Addr <= "0011011110010";
Trees_din <= "00000000000000000001001000010000";
wait for Clk_period;
Addr <= "0011011110011";
Trees_din <= "00000001000000000100000100001000";
wait for Clk_period;
Addr <= "0011011110100";
Trees_din <= "00000011000000000100101100000100";
wait for Clk_period;
Addr <= "0011011110101";
Trees_din <= "00000000001000100001110010111101";
wait for Clk_period;
Addr <= "0011011110110";
Trees_din <= "00000000000011010001110010111101";
wait for Clk_period;
Addr <= "0011011110111";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "0011011111000";
Trees_din <= "00000000000000100001110010111101";
wait for Clk_period;
Addr <= "0011011111001";
Trees_din <= "00000000010010100001110010111101";
wait for Clk_period;
Addr <= "0011011111010";
Trees_din <= "00000010000000000000100100001000";
wait for Clk_period;
Addr <= "0011011111011";
Trees_din <= "00000001000000000101011000000100";
wait for Clk_period;
Addr <= "0011011111100";
Trees_din <= "00000000010010100001110010111101";
wait for Clk_period;
Addr <= "0011011111101";
Trees_din <= "00000000010111010001110010111101";
wait for Clk_period;
Addr <= "0011011111110";
Trees_din <= "00000101000000000011110100000100";
wait for Clk_period;
Addr <= "0011011111111";
Trees_din <= "00000000010100010001110010111101";
wait for Clk_period;
Addr <= "0011100000000";
Trees_din <= "00000000000001010001110010111101";
wait for Clk_period;
Addr <= "0011100000001";
Trees_din <= "00000110000000000001110100010000";
wait for Clk_period;
Addr <= "0011100000010";
Trees_din <= "00000010000000000100011100001000";
wait for Clk_period;
Addr <= "0011100000011";
Trees_din <= "00000000000000000000111100000100";
wait for Clk_period;
Addr <= "0011100000100";
Trees_din <= "00000000001110010001110010111101";
wait for Clk_period;
Addr <= "0011100000101";
Trees_din <= "00000000000001000001110010111101";
wait for Clk_period;
Addr <= "0011100000110";
Trees_din <= "00000000000000000011111000000100";
wait for Clk_period;
Addr <= "0011100000111";
Trees_din <= "00000000010010110001110010111101";
wait for Clk_period;
Addr <= "0011100001000";
Trees_din <= "00000000001010000001110010111101";
wait for Clk_period;
Addr <= "0011100001001";
Trees_din <= "00000001000000000011111000001000";
wait for Clk_period;
Addr <= "0011100001010";
Trees_din <= "00000010000000000100101000000100";
wait for Clk_period;
Addr <= "0011100001011";
Trees_din <= "00000000010111000001110010111101";
wait for Clk_period;
Addr <= "0011100001100";
Trees_din <= "00000000010100110001110010111101";
wait for Clk_period;
Addr <= "0011100001101";
Trees_din <= "00000101000000000101111000000100";
wait for Clk_period;
Addr <= "0011100001110";
Trees_din <= "00000000000100110001110010111101";
wait for Clk_period;
Addr <= "0011100001111";
Trees_din <= "00000000010101100001110010111101";
wait for Clk_period;
Addr <= "0011100010000";
Trees_din <= "00000100000000000001010000100000";
wait for Clk_period;
Addr <= "0011100010001";
Trees_din <= "00000001000000000000001000010000";
wait for Clk_period;
Addr <= "0011100010010";
Trees_din <= "00000101000000000011001100001000";
wait for Clk_period;
Addr <= "0011100010011";
Trees_din <= "00000011000000000010011100000100";
wait for Clk_period;
Addr <= "0011100010100";
Trees_din <= "00000000000111100001110010111101";
wait for Clk_period;
Addr <= "0011100010101";
Trees_din <= "00000000001000000001110010111101";
wait for Clk_period;
Addr <= "0011100010110";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "0011100010111";
Trees_din <= "00000000010010000001110010111101";
wait for Clk_period;
Addr <= "0011100011000";
Trees_din <= "00000000010100100001110010111101";
wait for Clk_period;
Addr <= "0011100011001";
Trees_din <= "00000100000000000100110000001000";
wait for Clk_period;
Addr <= "0011100011010";
Trees_din <= "00000110000000000001101100000100";
wait for Clk_period;
Addr <= "0011100011011";
Trees_din <= "00000000010101010001110010111101";
wait for Clk_period;
Addr <= "0011100011100";
Trees_din <= "00000000000111110001110010111101";
wait for Clk_period;
Addr <= "0011100011101";
Trees_din <= "00000110000000000101111000000100";
wait for Clk_period;
Addr <= "0011100011110";
Trees_din <= "00000000010110000001110010111101";
wait for Clk_period;
Addr <= "0011100011111";
Trees_din <= "00000000000111010001110010111101";
wait for Clk_period;
Addr <= "0011100100000";
Trees_din <= "00000011000000000100011000010000";
wait for Clk_period;
Addr <= "0011100100001";
Trees_din <= "00000011000000000000010100001000";
wait for Clk_period;
Addr <= "0011100100010";
Trees_din <= "00000000000000000011100100000100";
wait for Clk_period;
Addr <= "0011100100011";
Trees_din <= "00000000000100110001110010111101";
wait for Clk_period;
Addr <= "0011100100100";
Trees_din <= "00000000001001010001110010111101";
wait for Clk_period;
Addr <= "0011100100101";
Trees_din <= "00000011000000000011000000000100";
wait for Clk_period;
Addr <= "0011100100110";
Trees_din <= "00000000010001000001110010111101";
wait for Clk_period;
Addr <= "0011100100111";
Trees_din <= "00000000000101000001110010111101";
wait for Clk_period;
Addr <= "0011100101000";
Trees_din <= "00000010000000000000000100001000";
wait for Clk_period;
Addr <= "0011100101001";
Trees_din <= "00000000000000000100101000000100";
wait for Clk_period;
Addr <= "0011100101010";
Trees_din <= "00000000001001010001110010111101";
wait for Clk_period;
Addr <= "0011100101011";
Trees_din <= "00000000001101100001110010111101";
wait for Clk_period;
Addr <= "0011100101100";
Trees_din <= "00000100000000000010010100000100";
wait for Clk_period;
Addr <= "0011100101101";
Trees_din <= "00000000010110100001110010111101";
wait for Clk_period;
Addr <= "0011100101110";
Trees_din <= "00000000000001110001110010111101";
wait for Clk_period;



----------tree 14-------------------

Addr <= "0011100101111";
Trees_din <= "00000001000000000100000110000000";
wait for Clk_period;
Addr <= "0011100110000";
Trees_din <= "00000010000000000100110101000000";
wait for Clk_period;
Addr <= "0011100110001";
Trees_din <= "00000010000000000100011100100000";
wait for Clk_period;
Addr <= "0011100110010";
Trees_din <= "00000001000000000010011100010000";
wait for Clk_period;
Addr <= "0011100110011";
Trees_din <= "00000100000000000110001000001000";
wait for Clk_period;
Addr <= "0011100110100";
Trees_din <= "00000110000000000011101100000100";
wait for Clk_period;
Addr <= "0011100110101";
Trees_din <= "00000000000101000001111010111011";
wait for Clk_period;
Addr <= "0011100110110";
Trees_din <= "00000000000000010001111010111011";
wait for Clk_period;
Addr <= "0011100110111";
Trees_din <= "00000011000000000100001000000100";
wait for Clk_period;
Addr <= "0011100111000";
Trees_din <= "00000000001110100001111010111011";
wait for Clk_period;
Addr <= "0011100111001";
Trees_din <= "00000000001110100001111010111011";
wait for Clk_period;
Addr <= "0011100111010";
Trees_din <= "00000101000000000010011000001000";
wait for Clk_period;
Addr <= "0011100111011";
Trees_din <= "00000110000000000011110100000100";
wait for Clk_period;
Addr <= "0011100111100";
Trees_din <= "00000000001010010001111010111011";
wait for Clk_period;
Addr <= "0011100111101";
Trees_din <= "00000000010011110001111010111011";
wait for Clk_period;
Addr <= "0011100111110";
Trees_din <= "00000111000000000000110000000100";
wait for Clk_period;
Addr <= "0011100111111";
Trees_din <= "00000000000011010001111010111011";
wait for Clk_period;
Addr <= "0011101000000";
Trees_din <= "00000000010101000001111010111011";
wait for Clk_period;
Addr <= "0011101000001";
Trees_din <= "00000000000000000011010000010000";
wait for Clk_period;
Addr <= "0011101000010";
Trees_din <= "00000000000000000100011100001000";
wait for Clk_period;
Addr <= "0011101000011";
Trees_din <= "00000011000000000010011100000100";
wait for Clk_period;
Addr <= "0011101000100";
Trees_din <= "00000000000101100001111010111011";
wait for Clk_period;
Addr <= "0011101000101";
Trees_din <= "00000000000011010001111010111011";
wait for Clk_period;
Addr <= "0011101000110";
Trees_din <= "00000001000000000011000000000100";
wait for Clk_period;
Addr <= "0011101000111";
Trees_din <= "00000000000011110001111010111011";
wait for Clk_period;
Addr <= "0011101001000";
Trees_din <= "00000000000011110001111010111011";
wait for Clk_period;
Addr <= "0011101001001";
Trees_din <= "00000110000000000010001000001000";
wait for Clk_period;
Addr <= "0011101001010";
Trees_din <= "00000110000000000000111100000100";
wait for Clk_period;
Addr <= "0011101001011";
Trees_din <= "00000000001001010001111010111011";
wait for Clk_period;
Addr <= "0011101001100";
Trees_din <= "00000000001100010001111010111011";
wait for Clk_period;
Addr <= "0011101001101";
Trees_din <= "00000101000000000001100100000100";
wait for Clk_period;
Addr <= "0011101001110";
Trees_din <= "00000000010101110001111010111011";
wait for Clk_period;
Addr <= "0011101001111";
Trees_din <= "00000000000011000001111010111011";
wait for Clk_period;
Addr <= "0011101010000";
Trees_din <= "00000001000000000010000100100000";
wait for Clk_period;
Addr <= "0011101010001";
Trees_din <= "00000000000000000000100000010000";
wait for Clk_period;
Addr <= "0011101010010";
Trees_din <= "00000110000000000000000100001000";
wait for Clk_period;
Addr <= "0011101010011";
Trees_din <= "00000110000000000001110000000100";
wait for Clk_period;
Addr <= "0011101010100";
Trees_din <= "00000000001100110001111010111011";
wait for Clk_period;
Addr <= "0011101010101";
Trees_din <= "00000000001010110001111010111011";
wait for Clk_period;
Addr <= "0011101010110";
Trees_din <= "00000000000000000101101000000100";
wait for Clk_period;
Addr <= "0011101010111";
Trees_din <= "00000000001111010001111010111011";
wait for Clk_period;
Addr <= "0011101011000";
Trees_din <= "00000000001001110001111010111011";
wait for Clk_period;
Addr <= "0011101011001";
Trees_din <= "00000000000000000101110100001000";
wait for Clk_period;
Addr <= "0011101011010";
Trees_din <= "00000110000000000011110000000100";
wait for Clk_period;
Addr <= "0011101011011";
Trees_din <= "00000000000110110001111010111011";
wait for Clk_period;
Addr <= "0011101011100";
Trees_din <= "00000000010100100001111010111011";
wait for Clk_period;
Addr <= "0011101011101";
Trees_din <= "00000010000000000000100000000100";
wait for Clk_period;
Addr <= "0011101011110";
Trees_din <= "00000000000000110001111010111011";
wait for Clk_period;
Addr <= "0011101011111";
Trees_din <= "00000000010100010001111010111011";
wait for Clk_period;
Addr <= "0011101100000";
Trees_din <= "00000111000000000010001100010000";
wait for Clk_period;
Addr <= "0011101100001";
Trees_din <= "00000001000000000010010100001000";
wait for Clk_period;
Addr <= "0011101100010";
Trees_din <= "00000001000000000101100100000100";
wait for Clk_period;
Addr <= "0011101100011";
Trees_din <= "00000000001011110001111010111011";
wait for Clk_period;
Addr <= "0011101100100";
Trees_din <= "00000000010000010001111010111011";
wait for Clk_period;
Addr <= "0011101100101";
Trees_din <= "00000101000000000110001000000100";
wait for Clk_period;
Addr <= "0011101100110";
Trees_din <= "00000000001101010001111010111011";
wait for Clk_period;
Addr <= "0011101100111";
Trees_din <= "00000000011000100001111010111011";
wait for Clk_period;
Addr <= "0011101101000";
Trees_din <= "00000001000000000101011000001000";
wait for Clk_period;
Addr <= "0011101101001";
Trees_din <= "00000110000000000010110100000100";
wait for Clk_period;
Addr <= "0011101101010";
Trees_din <= "00000000001011010001111010111011";
wait for Clk_period;
Addr <= "0011101101011";
Trees_din <= "00000000000010000001111010111011";
wait for Clk_period;
Addr <= "0011101101100";
Trees_din <= "00000110000000000000100000000100";
wait for Clk_period;
Addr <= "0011101101101";
Trees_din <= "00000000011001000001111010111011";
wait for Clk_period;
Addr <= "0011101101110";
Trees_din <= "00000000010111000001111010111011";
wait for Clk_period;
Addr <= "0011101101111";
Trees_din <= "00000000000000000010011101000000";
wait for Clk_period;
Addr <= "0011101110000";
Trees_din <= "00000001000000000101101100100000";
wait for Clk_period;
Addr <= "0011101110001";
Trees_din <= "00000100000000000001101100010000";
wait for Clk_period;
Addr <= "0011101110010";
Trees_din <= "00000000000000000010111100001000";
wait for Clk_period;
Addr <= "0011101110011";
Trees_din <= "00000011000000000100101100000100";
wait for Clk_period;
Addr <= "0011101110100";
Trees_din <= "00000000000010010001111010111011";
wait for Clk_period;
Addr <= "0011101110101";
Trees_din <= "00000000001100010001111010111011";
wait for Clk_period;
Addr <= "0011101110110";
Trees_din <= "00000100000000000000101100000100";
wait for Clk_period;
Addr <= "0011101110111";
Trees_din <= "00000000000011100001111010111011";
wait for Clk_period;
Addr <= "0011101111000";
Trees_din <= "00000000001110100001111010111011";
wait for Clk_period;
Addr <= "0011101111001";
Trees_din <= "00000100000000000101100000001000";
wait for Clk_period;
Addr <= "0011101111010";
Trees_din <= "00000010000000000110000000000100";
wait for Clk_period;
Addr <= "0011101111011";
Trees_din <= "00000000010010000001111010111011";
wait for Clk_period;
Addr <= "0011101111100";
Trees_din <= "00000000000110100001111010111011";
wait for Clk_period;
Addr <= "0011101111101";
Trees_din <= "00000101000000000101001000000100";
wait for Clk_period;
Addr <= "0011101111110";
Trees_din <= "00000000010010000001111010111011";
wait for Clk_period;
Addr <= "0011101111111";
Trees_din <= "00000000010011100001111010111011";
wait for Clk_period;
Addr <= "0011110000000";
Trees_din <= "00000111000000000000000100010000";
wait for Clk_period;
Addr <= "0011110000001";
Trees_din <= "00000101000000000001010100001000";
wait for Clk_period;
Addr <= "0011110000010";
Trees_din <= "00000101000000000101010000000100";
wait for Clk_period;
Addr <= "0011110000011";
Trees_din <= "00000000000011100001111010111011";
wait for Clk_period;
Addr <= "0011110000100";
Trees_din <= "00000000010011100001111010111011";
wait for Clk_period;
Addr <= "0011110000101";
Trees_din <= "00000010000000000100001100000100";
wait for Clk_period;
Addr <= "0011110000110";
Trees_din <= "00000000001100110001111010111011";
wait for Clk_period;
Addr <= "0011110000111";
Trees_din <= "00000000000010110001111010111011";
wait for Clk_period;
Addr <= "0011110001000";
Trees_din <= "00000010000000000000101000001000";
wait for Clk_period;
Addr <= "0011110001001";
Trees_din <= "00000100000000000000001100000100";
wait for Clk_period;
Addr <= "0011110001010";
Trees_din <= "00000000000001110001111010111011";
wait for Clk_period;
Addr <= "0011110001011";
Trees_din <= "00000000010011100001111010111011";
wait for Clk_period;
Addr <= "0011110001100";
Trees_din <= "00000011000000000001101000000100";
wait for Clk_period;
Addr <= "0011110001101";
Trees_din <= "00000000000111000001111010111011";
wait for Clk_period;
Addr <= "0011110001110";
Trees_din <= "00000000011000110001111010111011";
wait for Clk_period;
Addr <= "0011110001111";
Trees_din <= "00000101000000000101011000100000";
wait for Clk_period;
Addr <= "0011110010000";
Trees_din <= "00000111000000000010010100010000";
wait for Clk_period;
Addr <= "0011110010001";
Trees_din <= "00000111000000000100011000001000";
wait for Clk_period;
Addr <= "0011110010010";
Trees_din <= "00000001000000000000101100000100";
wait for Clk_period;
Addr <= "0011110010011";
Trees_din <= "00000000010010100001111010111011";
wait for Clk_period;
Addr <= "0011110010100";
Trees_din <= "00000000000110100001111010111011";
wait for Clk_period;
Addr <= "0011110010101";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "0011110010110";
Trees_din <= "00000000000010000001111010111011";
wait for Clk_period;
Addr <= "0011110010111";
Trees_din <= "00000000001110110001111010111011";
wait for Clk_period;
Addr <= "0011110011000";
Trees_din <= "00000101000000000001001000001000";
wait for Clk_period;
Addr <= "0011110011001";
Trees_din <= "00000000000000000100101100000100";
wait for Clk_period;
Addr <= "0011110011010";
Trees_din <= "00000000010100110001111010111011";
wait for Clk_period;
Addr <= "0011110011011";
Trees_din <= "00000000000010000001111010111011";
wait for Clk_period;
Addr <= "0011110011100";
Trees_din <= "00000011000000000101011000000100";
wait for Clk_period;
Addr <= "0011110011101";
Trees_din <= "00000000001100000001111010111011";
wait for Clk_period;
Addr <= "0011110011110";
Trees_din <= "00000000010011000001111010111011";
wait for Clk_period;
Addr <= "0011110011111";
Trees_din <= "00000000000000000001001100010000";
wait for Clk_period;
Addr <= "0011110100000";
Trees_din <= "00000110000000000101010000001000";
wait for Clk_period;
Addr <= "0011110100001";
Trees_din <= "00000001000000000011111000000100";
wait for Clk_period;
Addr <= "0011110100010";
Trees_din <= "00000000010010010001111010111011";
wait for Clk_period;
Addr <= "0011110100011";
Trees_din <= "00000000001101100001111010111011";
wait for Clk_period;
Addr <= "0011110100100";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "0011110100101";
Trees_din <= "00000000000100000001111010111011";
wait for Clk_period;
Addr <= "0011110100110";
Trees_din <= "00000000010111100001111010111011";
wait for Clk_period;
Addr <= "0011110100111";
Trees_din <= "00000101000000000011111000001000";
wait for Clk_period;
Addr <= "0011110101000";
Trees_din <= "00000010000000000010001000000100";
wait for Clk_period;
Addr <= "0011110101001";
Trees_din <= "00000000011000100001111010111011";
wait for Clk_period;
Addr <= "0011110101010";
Trees_din <= "00000000010010000001111010111011";
wait for Clk_period;
Addr <= "0011110101011";
Trees_din <= "00000010000000000101010000000100";
wait for Clk_period;
Addr <= "0011110101100";
Trees_din <= "00000000000111110001111010111011";
wait for Clk_period;
Addr <= "0011110101101";
Trees_din <= "00000000000110100001111010111011";
wait for Clk_period;



----------tree 15-------------------

Addr <= "0011110101110";
Trees_din <= "00000111000000000011010110000000";
wait for Clk_period;
Addr <= "0011110101111";
Trees_din <= "00000000000000000101101001000000";
wait for Clk_period;
Addr <= "0011110110000";
Trees_din <= "00000100000000000001010100100000";
wait for Clk_period;
Addr <= "0011110110001";
Trees_din <= "00000001000000000110000100010000";
wait for Clk_period;
Addr <= "0011110110010";
Trees_din <= "00000000000000000100110100001000";
wait for Clk_period;
Addr <= "0011110110011";
Trees_din <= "00000001000000000010110000000100";
wait for Clk_period;
Addr <= "0011110110100";
Trees_din <= "00000000010110110010000010110101";
wait for Clk_period;
Addr <= "0011110110101";
Trees_din <= "00000000001110100010000010110101";
wait for Clk_period;
Addr <= "0011110110110";
Trees_din <= "00000100000000000011100000000100";
wait for Clk_period;
Addr <= "0011110110111";
Trees_din <= "00000000011000110010000010110101";
wait for Clk_period;
Addr <= "0011110111000";
Trees_din <= "00000000000100000010000010110101";
wait for Clk_period;
Addr <= "0011110111001";
Trees_din <= "00000111000000000001110100001000";
wait for Clk_period;
Addr <= "0011110111010";
Trees_din <= "00000110000000000100010100000100";
wait for Clk_period;
Addr <= "0011110111011";
Trees_din <= "00000000001011010010000010110101";
wait for Clk_period;
Addr <= "0011110111100";
Trees_din <= "00000000000010010010000010110101";
wait for Clk_period;
Addr <= "0011110111101";
Trees_din <= "00000101000000000011001100000100";
wait for Clk_period;
Addr <= "0011110111110";
Trees_din <= "00000000000101010010000010110101";
wait for Clk_period;
Addr <= "0011110111111";
Trees_din <= "00000000000111110010000010110101";
wait for Clk_period;
Addr <= "0011111000000";
Trees_din <= "00000001000000000100010000010000";
wait for Clk_period;
Addr <= "0011111000001";
Trees_din <= "00000011000000000000011000001000";
wait for Clk_period;
Addr <= "0011111000010";
Trees_din <= "00000111000000000100101100000100";
wait for Clk_period;
Addr <= "0011111000011";
Trees_din <= "00000000011000010010000010110101";
wait for Clk_period;
Addr <= "0011111000100";
Trees_din <= "00000000010000010010000010110101";
wait for Clk_period;
Addr <= "0011111000101";
Trees_din <= "00000010000000000011011000000100";
wait for Clk_period;
Addr <= "0011111000110";
Trees_din <= "00000000010010110010000010110101";
wait for Clk_period;
Addr <= "0011111000111";
Trees_din <= "00000000000001100010000010110101";
wait for Clk_period;
Addr <= "0011111001000";
Trees_din <= "00000001000000000000011000001000";
wait for Clk_period;
Addr <= "0011111001001";
Trees_din <= "00000101000000000000100100000100";
wait for Clk_period;
Addr <= "0011111001010";
Trees_din <= "00000000010010100010000010110101";
wait for Clk_period;
Addr <= "0011111001011";
Trees_din <= "00000000000000110010000010110101";
wait for Clk_period;
Addr <= "0011111001100";
Trees_din <= "00000111000000000110001000000100";
wait for Clk_period;
Addr <= "0011111001101";
Trees_din <= "00000000000101000010000010110101";
wait for Clk_period;
Addr <= "0011111001110";
Trees_din <= "00000000000110000010000010110101";
wait for Clk_period;
Addr <= "0011111001111";
Trees_din <= "00000000000000000101110100100000";
wait for Clk_period;
Addr <= "0011111010000";
Trees_din <= "00000000000000000011001100010000";
wait for Clk_period;
Addr <= "0011111010001";
Trees_din <= "00000111000000000010001000001000";
wait for Clk_period;
Addr <= "0011111010010";
Trees_din <= "00000000000000000010110100000100";
wait for Clk_period;
Addr <= "0011111010011";
Trees_din <= "00000000000010100010000010110101";
wait for Clk_period;
Addr <= "0011111010100";
Trees_din <= "00000000001110100010000010110101";
wait for Clk_period;
Addr <= "0011111010101";
Trees_din <= "00000001000000000101110000000100";
wait for Clk_period;
Addr <= "0011111010110";
Trees_din <= "00000000000001100010000010110101";
wait for Clk_period;
Addr <= "0011111010111";
Trees_din <= "00000000001111100010000010110101";
wait for Clk_period;
Addr <= "0011111011000";
Trees_din <= "00000000000000000100101000001000";
wait for Clk_period;
Addr <= "0011111011001";
Trees_din <= "00000000000000000011011000000100";
wait for Clk_period;
Addr <= "0011111011010";
Trees_din <= "00000000010101000010000010110101";
wait for Clk_period;
Addr <= "0011111011011";
Trees_din <= "00000000000111010010000010110101";
wait for Clk_period;
Addr <= "0011111011100";
Trees_din <= "00000111000000000000010000000100";
wait for Clk_period;
Addr <= "0011111011101";
Trees_din <= "00000000000111100010000010110101";
wait for Clk_period;
Addr <= "0011111011110";
Trees_din <= "00000000000000010010000010110101";
wait for Clk_period;
Addr <= "0011111011111";
Trees_din <= "00000011000000000001010100010000";
wait for Clk_period;
Addr <= "0011111100000";
Trees_din <= "00000100000000000000100100001000";
wait for Clk_period;
Addr <= "0011111100001";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "0011111100010";
Trees_din <= "00000000001100110010000010110101";
wait for Clk_period;
Addr <= "0011111100011";
Trees_din <= "00000000001001100010000010110101";
wait for Clk_period;
Addr <= "0011111100100";
Trees_din <= "00000111000000000101111100000100";
wait for Clk_period;
Addr <= "0011111100101";
Trees_din <= "00000000001001100010000010110101";
wait for Clk_period;
Addr <= "0011111100110";
Trees_din <= "00000000001111110010000010110101";
wait for Clk_period;
Addr <= "0011111100111";
Trees_din <= "00000010000000000001110000001000";
wait for Clk_period;
Addr <= "0011111101000";
Trees_din <= "00000000000000000101111000000100";
wait for Clk_period;
Addr <= "0011111101001";
Trees_din <= "00000000010011010010000010110101";
wait for Clk_period;
Addr <= "0011111101010";
Trees_din <= "00000000010011010010000010110101";
wait for Clk_period;
Addr <= "0011111101011";
Trees_din <= "00000110000000000100000100000100";
wait for Clk_period;
Addr <= "0011111101100";
Trees_din <= "00000000000000100010000010110101";
wait for Clk_period;
Addr <= "0011111101101";
Trees_din <= "00000000001001110010000010110101";
wait for Clk_period;
Addr <= "0011111101110";
Trees_din <= "00000010000000000101100101000000";
wait for Clk_period;
Addr <= "0011111101111";
Trees_din <= "00000110000000000000000100100000";
wait for Clk_period;
Addr <= "0011111110000";
Trees_din <= "00000000000000000101001000010000";
wait for Clk_period;
Addr <= "0011111110001";
Trees_din <= "00000101000000000010110100001000";
wait for Clk_period;
Addr <= "0011111110010";
Trees_din <= "00000001000000000101010000000100";
wait for Clk_period;
Addr <= "0011111110011";
Trees_din <= "00000000010000110010000010110101";
wait for Clk_period;
Addr <= "0011111110100";
Trees_din <= "00000000010100000010000010110101";
wait for Clk_period;
Addr <= "0011111110101";
Trees_din <= "00000101000000000010101100000100";
wait for Clk_period;
Addr <= "0011111110110";
Trees_din <= "00000000001111010010000010110101";
wait for Clk_period;
Addr <= "0011111110111";
Trees_din <= "00000000001011110010000010110101";
wait for Clk_period;
Addr <= "0011111111000";
Trees_din <= "00000010000000000100101100001000";
wait for Clk_period;
Addr <= "0011111111001";
Trees_din <= "00000001000000000100100100000100";
wait for Clk_period;
Addr <= "0011111111010";
Trees_din <= "00000000001010010010000010110101";
wait for Clk_period;
Addr <= "0011111111011";
Trees_din <= "00000000000100000010000010110101";
wait for Clk_period;
Addr <= "0011111111100";
Trees_din <= "00000000000000000010010000000100";
wait for Clk_period;
Addr <= "0011111111101";
Trees_din <= "00000000001100100010000010110101";
wait for Clk_period;
Addr <= "0011111111110";
Trees_din <= "00000000010111000010000010110101";
wait for Clk_period;
Addr <= "0011111111111";
Trees_din <= "00000010000000000101101000010000";
wait for Clk_period;
Addr <= "0100000000000";
Trees_din <= "00000000000000000101001000001000";
wait for Clk_period;
Addr <= "0100000000001";
Trees_din <= "00000110000000000101010000000100";
wait for Clk_period;
Addr <= "0100000000010";
Trees_din <= "00000000001100110010000010110101";
wait for Clk_period;
Addr <= "0100000000011";
Trees_din <= "00000000000001010010000010110101";
wait for Clk_period;
Addr <= "0100000000100";
Trees_din <= "00000110000000000100111100000100";
wait for Clk_period;
Addr <= "0100000000101";
Trees_din <= "00000000010001110010000010110101";
wait for Clk_period;
Addr <= "0100000000110";
Trees_din <= "00000000001110010010000010110101";
wait for Clk_period;
Addr <= "0100000000111";
Trees_din <= "00000010000000000000101000001000";
wait for Clk_period;
Addr <= "0100000001000";
Trees_din <= "00000011000000000001111000000100";
wait for Clk_period;
Addr <= "0100000001001";
Trees_din <= "00000000000101100010000010110101";
wait for Clk_period;
Addr <= "0100000001010";
Trees_din <= "00000000010101010010000010110101";
wait for Clk_period;
Addr <= "0100000001011";
Trees_din <= "00000110000000000101011100000100";
wait for Clk_period;
Addr <= "0100000001100";
Trees_din <= "00000000000101000010000010110101";
wait for Clk_period;
Addr <= "0100000001101";
Trees_din <= "00000000001110010010000010110101";
wait for Clk_period;
Addr <= "0100000001110";
Trees_din <= "00000110000000000101100100100000";
wait for Clk_period;
Addr <= "0100000001111";
Trees_din <= "00000010000000000100010100010000";
wait for Clk_period;
Addr <= "0100000010000";
Trees_din <= "00000010000000000011100100001000";
wait for Clk_period;
Addr <= "0100000010001";
Trees_din <= "00000001000000000000111100000100";
wait for Clk_period;
Addr <= "0100000010010";
Trees_din <= "00000000010101010010000010110101";
wait for Clk_period;
Addr <= "0100000010011";
Trees_din <= "00000000001100100010000010110101";
wait for Clk_period;
Addr <= "0100000010100";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "0100000010101";
Trees_din <= "00000000010110000010000010110101";
wait for Clk_period;
Addr <= "0100000010110";
Trees_din <= "00000000010001100010000010110101";
wait for Clk_period;
Addr <= "0100000010111";
Trees_din <= "00000100000000000001001100001000";
wait for Clk_period;
Addr <= "0100000011000";
Trees_din <= "00000101000000000110000100000100";
wait for Clk_period;
Addr <= "0100000011001";
Trees_din <= "00000000001011100010000010110101";
wait for Clk_period;
Addr <= "0100000011010";
Trees_din <= "00000000000000000010000010110101";
wait for Clk_period;
Addr <= "0100000011011";
Trees_din <= "00000001000000000001011000000100";
wait for Clk_period;
Addr <= "0100000011100";
Trees_din <= "00000000010111110010000010110101";
wait for Clk_period;
Addr <= "0100000011101";
Trees_din <= "00000000001001000010000010110101";
wait for Clk_period;
Addr <= "0100000011110";
Trees_din <= "00000101000000000010001100010000";
wait for Clk_period;
Addr <= "0100000011111";
Trees_din <= "00000001000000000001011000001000";
wait for Clk_period;
Addr <= "0100000100000";
Trees_din <= "00000100000000000010010100000100";
wait for Clk_period;
Addr <= "0100000100001";
Trees_din <= "00000000011001000010000010110101";
wait for Clk_period;
Addr <= "0100000100010";
Trees_din <= "00000000001011000010000010110101";
wait for Clk_period;
Addr <= "0100000100011";
Trees_din <= "00000011000000000000111000000100";
wait for Clk_period;
Addr <= "0100000100100";
Trees_din <= "00000000010011110010000010110101";
wait for Clk_period;
Addr <= "0100000100101";
Trees_din <= "00000000001010100010000010110101";
wait for Clk_period;
Addr <= "0100000100110";
Trees_din <= "00000110000000000010011100001000";
wait for Clk_period;
Addr <= "0100000100111";
Trees_din <= "00000001000000000101000100000100";
wait for Clk_period;
Addr <= "0100000101000";
Trees_din <= "00000000010110100010000010110101";
wait for Clk_period;
Addr <= "0100000101001";
Trees_din <= "00000000010000100010000010110101";
wait for Clk_period;
Addr <= "0100000101010";
Trees_din <= "00000100000000000010011100000100";
wait for Clk_period;
Addr <= "0100000101011";
Trees_din <= "00000000000000110010000010110101";
wait for Clk_period;
Addr <= "0100000101100";
Trees_din <= "00000000000010100010000010110101";
wait for Clk_period;



----------tree 16-------------------

Addr <= "0100000101101";
Trees_din <= "00000100000000000000110010000000";
wait for Clk_period;
Addr <= "0100000101110";
Trees_din <= "00000001000000000001011101000000";
wait for Clk_period;
Addr <= "0100000101111";
Trees_din <= "00000010000000000101111000100000";
wait for Clk_period;
Addr <= "0100000110000";
Trees_din <= "00000011000000000001011000010000";
wait for Clk_period;
Addr <= "0100000110001";
Trees_din <= "00000011000000000101100100001000";
wait for Clk_period;
Addr <= "0100000110010";
Trees_din <= "00000101000000000101111000000100";
wait for Clk_period;
Addr <= "0100000110011";
Trees_din <= "00000000000110010010001010110001";
wait for Clk_period;
Addr <= "0100000110100";
Trees_din <= "00000000001110110010001010110001";
wait for Clk_period;
Addr <= "0100000110101";
Trees_din <= "00000110000000000001101000000100";
wait for Clk_period;
Addr <= "0100000110110";
Trees_din <= "00000000001101110010001010110001";
wait for Clk_period;
Addr <= "0100000110111";
Trees_din <= "00000000000100110010001010110001";
wait for Clk_period;
Addr <= "0100000111000";
Trees_din <= "00000001000000000001000100001000";
wait for Clk_period;
Addr <= "0100000111001";
Trees_din <= "00000010000000000000001100000100";
wait for Clk_period;
Addr <= "0100000111010";
Trees_din <= "00000000001010010010001010110001";
wait for Clk_period;
Addr <= "0100000111011";
Trees_din <= "00000000001101000010001010110001";
wait for Clk_period;
Addr <= "0100000111100";
Trees_din <= "00000110000000000001001000000100";
wait for Clk_period;
Addr <= "0100000111101";
Trees_din <= "00000000000000010010001010110001";
wait for Clk_period;
Addr <= "0100000111110";
Trees_din <= "00000000000000110010001010110001";
wait for Clk_period;
Addr <= "0100000111111";
Trees_din <= "00000110000000000100101000010000";
wait for Clk_period;
Addr <= "0100001000000";
Trees_din <= "00000111000000000011100000001000";
wait for Clk_period;
Addr <= "0100001000001";
Trees_din <= "00000111000000000011111000000100";
wait for Clk_period;
Addr <= "0100001000010";
Trees_din <= "00000000001110100010001010110001";
wait for Clk_period;
Addr <= "0100001000011";
Trees_din <= "00000000000100110010001010110001";
wait for Clk_period;
Addr <= "0100001000100";
Trees_din <= "00000001000000000000000100000100";
wait for Clk_period;
Addr <= "0100001000101";
Trees_din <= "00000000001000110010001010110001";
wait for Clk_period;
Addr <= "0100001000110";
Trees_din <= "00000000001100000010001010110001";
wait for Clk_period;
Addr <= "0100001000111";
Trees_din <= "00000000000000000100101100001000";
wait for Clk_period;
Addr <= "0100001001000";
Trees_din <= "00000110000000000010010000000100";
wait for Clk_period;
Addr <= "0100001001001";
Trees_din <= "00000000000010010010001010110001";
wait for Clk_period;
Addr <= "0100001001010";
Trees_din <= "00000000010001000010001010110001";
wait for Clk_period;
Addr <= "0100001001011";
Trees_din <= "00000000000000000110001000000100";
wait for Clk_period;
Addr <= "0100001001100";
Trees_din <= "00000000000011100010001010110001";
wait for Clk_period;
Addr <= "0100001001101";
Trees_din <= "00000000010000110010001010110001";
wait for Clk_period;
Addr <= "0100001001110";
Trees_din <= "00000011000000000100000000100000";
wait for Clk_period;
Addr <= "0100001001111";
Trees_din <= "00000100000000000000100000010000";
wait for Clk_period;
Addr <= "0100001010000";
Trees_din <= "00000011000000000100111100001000";
wait for Clk_period;
Addr <= "0100001010001";
Trees_din <= "00000110000000000100010100000100";
wait for Clk_period;
Addr <= "0100001010010";
Trees_din <= "00000000001100100010001010110001";
wait for Clk_period;
Addr <= "0100001010011";
Trees_din <= "00000000001011110010001010110001";
wait for Clk_period;
Addr <= "0100001010100";
Trees_din <= "00000111000000000100000100000100";
wait for Clk_period;
Addr <= "0100001010101";
Trees_din <= "00000000001100000010001010110001";
wait for Clk_period;
Addr <= "0100001010110";
Trees_din <= "00000000001010000010001010110001";
wait for Clk_period;
Addr <= "0100001010111";
Trees_din <= "00000001000000000010001100001000";
wait for Clk_period;
Addr <= "0100001011000";
Trees_din <= "00000010000000000101010000000100";
wait for Clk_period;
Addr <= "0100001011001";
Trees_din <= "00000000010011000010001010110001";
wait for Clk_period;
Addr <= "0100001011010";
Trees_din <= "00000000010111010010001010110001";
wait for Clk_period;
Addr <= "0100001011011";
Trees_din <= "00000100000000000011110000000100";
wait for Clk_period;
Addr <= "0100001011100";
Trees_din <= "00000000001011110010001010110001";
wait for Clk_period;
Addr <= "0100001011101";
Trees_din <= "00000000011000110010001010110001";
wait for Clk_period;
Addr <= "0100001011110";
Trees_din <= "00000100000000000000010000010000";
wait for Clk_period;
Addr <= "0100001011111";
Trees_din <= "00000100000000000010011000001000";
wait for Clk_period;
Addr <= "0100001100000";
Trees_din <= "00000100000000000100010000000100";
wait for Clk_period;
Addr <= "0100001100001";
Trees_din <= "00000000011000100010001010110001";
wait for Clk_period;
Addr <= "0100001100010";
Trees_din <= "00000000000101000010001010110001";
wait for Clk_period;
Addr <= "0100001100011";
Trees_din <= "00000010000000000010000100000100";
wait for Clk_period;
Addr <= "0100001100100";
Trees_din <= "00000000001111000010001010110001";
wait for Clk_period;
Addr <= "0100001100101";
Trees_din <= "00000000000000000010001010110001";
wait for Clk_period;
Addr <= "0100001100110";
Trees_din <= "00000001000000000001111100001000";
wait for Clk_period;
Addr <= "0100001100111";
Trees_din <= "00000101000000000011110000000100";
wait for Clk_period;
Addr <= "0100001101000";
Trees_din <= "00000000010011110010001010110001";
wait for Clk_period;
Addr <= "0100001101001";
Trees_din <= "00000000010000100010001010110001";
wait for Clk_period;
Addr <= "0100001101010";
Trees_din <= "00000001000000000001101000000100";
wait for Clk_period;
Addr <= "0100001101011";
Trees_din <= "00000000010110110010001010110001";
wait for Clk_period;
Addr <= "0100001101100";
Trees_din <= "00000000010100110010001010110001";
wait for Clk_period;
Addr <= "0100001101101";
Trees_din <= "00000101000000000101111001000000";
wait for Clk_period;
Addr <= "0100001101110";
Trees_din <= "00000110000000000010110000100000";
wait for Clk_period;
Addr <= "0100001101111";
Trees_din <= "00000011000000000100001000010000";
wait for Clk_period;
Addr <= "0100001110000";
Trees_din <= "00000110000000000001101100001000";
wait for Clk_period;
Addr <= "0100001110001";
Trees_din <= "00000000000000000000010000000100";
wait for Clk_period;
Addr <= "0100001110010";
Trees_din <= "00000000000110100010001010110001";
wait for Clk_period;
Addr <= "0100001110011";
Trees_din <= "00000000001101110010001010110001";
wait for Clk_period;
Addr <= "0100001110100";
Trees_din <= "00000111000000000001000100000100";
wait for Clk_period;
Addr <= "0100001110101";
Trees_din <= "00000000010001010010001010110001";
wait for Clk_period;
Addr <= "0100001110110";
Trees_din <= "00000000010110010010001010110001";
wait for Clk_period;
Addr <= "0100001110111";
Trees_din <= "00000101000000000000010000001000";
wait for Clk_period;
Addr <= "0100001111000";
Trees_din <= "00000001000000000101101100000100";
wait for Clk_period;
Addr <= "0100001111001";
Trees_din <= "00000000010010010010001010110001";
wait for Clk_period;
Addr <= "0100001111010";
Trees_din <= "00000000001000000010001010110001";
wait for Clk_period;
Addr <= "0100001111011";
Trees_din <= "00000110000000000110001100000100";
wait for Clk_period;
Addr <= "0100001111100";
Trees_din <= "00000000001101100010001010110001";
wait for Clk_period;
Addr <= "0100001111101";
Trees_din <= "00000000000000000010001010110001";
wait for Clk_period;
Addr <= "0100001111110";
Trees_din <= "00000010000000000010011000010000";
wait for Clk_period;
Addr <= "0100001111111";
Trees_din <= "00000111000000000101011000001000";
wait for Clk_period;
Addr <= "0100010000000";
Trees_din <= "00000111000000000011110100000100";
wait for Clk_period;
Addr <= "0100010000001";
Trees_din <= "00000000011001000010001010110001";
wait for Clk_period;
Addr <= "0100010000010";
Trees_din <= "00000000000111010010001010110001";
wait for Clk_period;
Addr <= "0100010000011";
Trees_din <= "00000001000000000011100100000100";
wait for Clk_period;
Addr <= "0100010000100";
Trees_din <= "00000000010111100010001010110001";
wait for Clk_period;
Addr <= "0100010000101";
Trees_din <= "00000000010000110010001010110001";
wait for Clk_period;
Addr <= "0100010000110";
Trees_din <= "00000110000000000100111000001000";
wait for Clk_period;
Addr <= "0100010000111";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "0100010001000";
Trees_din <= "00000000010110000010001010110001";
wait for Clk_period;
Addr <= "0100010001001";
Trees_din <= "00000000001011100010001010110001";
wait for Clk_period;
Addr <= "0100010001010";
Trees_din <= "00000110000000000011101100000100";
wait for Clk_period;
Addr <= "0100010001011";
Trees_din <= "00000000001111000010001010110001";
wait for Clk_period;
Addr <= "0100010001100";
Trees_din <= "00000000001101010010001010110001";
wait for Clk_period;
Addr <= "0100010001101";
Trees_din <= "00000011000000000011001000100000";
wait for Clk_period;
Addr <= "0100010001110";
Trees_din <= "00000111000000000011011000010000";
wait for Clk_period;
Addr <= "0100010001111";
Trees_din <= "00000111000000000001011000001000";
wait for Clk_period;
Addr <= "0100010010000";
Trees_din <= "00000111000000000110010000000100";
wait for Clk_period;
Addr <= "0100010010001";
Trees_din <= "00000000010101010010001010110001";
wait for Clk_period;
Addr <= "0100010010010";
Trees_din <= "00000000000001000010001010110001";
wait for Clk_period;
Addr <= "0100010010011";
Trees_din <= "00000110000000000100110100000100";
wait for Clk_period;
Addr <= "0100010010100";
Trees_din <= "00000000001111110010001010110001";
wait for Clk_period;
Addr <= "0100010010101";
Trees_din <= "00000000000111110010001010110001";
wait for Clk_period;
Addr <= "0100010010110";
Trees_din <= "00000100000000000000110000001000";
wait for Clk_period;
Addr <= "0100010010111";
Trees_din <= "00000001000000000001101100000100";
wait for Clk_period;
Addr <= "0100010011000";
Trees_din <= "00000000001001110010001010110001";
wait for Clk_period;
Addr <= "0100010011001";
Trees_din <= "00000000001001010010001010110001";
wait for Clk_period;
Addr <= "0100010011010";
Trees_din <= "00000111000000000000011000000100";
wait for Clk_period;
Addr <= "0100010011011";
Trees_din <= "00000000000101010010001010110001";
wait for Clk_period;
Addr <= "0100010011100";
Trees_din <= "00000000000100110010001010110001";
wait for Clk_period;
Addr <= "0100010011101";
Trees_din <= "00000111000000000101000100010000";
wait for Clk_period;
Addr <= "0100010011110";
Trees_din <= "00000001000000000000111100001000";
wait for Clk_period;
Addr <= "0100010011111";
Trees_din <= "00000100000000000100000100000100";
wait for Clk_period;
Addr <= "0100010100000";
Trees_din <= "00000000000001010010001010110001";
wait for Clk_period;
Addr <= "0100010100001";
Trees_din <= "00000000010011000010001010110001";
wait for Clk_period;
Addr <= "0100010100010";
Trees_din <= "00000001000000000001101100000100";
wait for Clk_period;
Addr <= "0100010100011";
Trees_din <= "00000000000100110010001010110001";
wait for Clk_period;
Addr <= "0100010100100";
Trees_din <= "00000000000101000010001010110001";
wait for Clk_period;
Addr <= "0100010100101";
Trees_din <= "00000110000000000100010100001000";
wait for Clk_period;
Addr <= "0100010100110";
Trees_din <= "00000011000000000101110000000100";
wait for Clk_period;
Addr <= "0100010100111";
Trees_din <= "00000000000011100010001010110001";
wait for Clk_period;
Addr <= "0100010101000";
Trees_din <= "00000000000010100010001010110001";
wait for Clk_period;
Addr <= "0100010101001";
Trees_din <= "00000001000000000101101000000100";
wait for Clk_period;
Addr <= "0100010101010";
Trees_din <= "00000000000101100010001010110001";
wait for Clk_period;
Addr <= "0100010101011";
Trees_din <= "00000000001000110010001010110001";
wait for Clk_period;



----------tree 17-------------------

Addr <= "0100010101100";
Trees_din <= "00000111000000000100111110000000";
wait for Clk_period;
Addr <= "0100010101101";
Trees_din <= "00000001000000000101110101000000";
wait for Clk_period;
Addr <= "0100010101110";
Trees_din <= "00000101000000000100101000100000";
wait for Clk_period;
Addr <= "0100010101111";
Trees_din <= "00000010000000000011010000010000";
wait for Clk_period;
Addr <= "0100010110000";
Trees_din <= "00000101000000000000101000001000";
wait for Clk_period;
Addr <= "0100010110001";
Trees_din <= "00000100000000000011011100000100";
wait for Clk_period;
Addr <= "0100010110010";
Trees_din <= "00000000010100000010010010101101";
wait for Clk_period;
Addr <= "0100010110011";
Trees_din <= "00000000000111100010010010101101";
wait for Clk_period;
Addr <= "0100010110100";
Trees_din <= "00000010000000000010011100000100";
wait for Clk_period;
Addr <= "0100010110101";
Trees_din <= "00000000010111010010010010101101";
wait for Clk_period;
Addr <= "0100010110110";
Trees_din <= "00000000000101100010010010101101";
wait for Clk_period;
Addr <= "0100010110111";
Trees_din <= "00000110000000000100010000001000";
wait for Clk_period;
Addr <= "0100010111000";
Trees_din <= "00000001000000000001110100000100";
wait for Clk_period;
Addr <= "0100010111001";
Trees_din <= "00000000001101010010010010101101";
wait for Clk_period;
Addr <= "0100010111010";
Trees_din <= "00000000000111010010010010101101";
wait for Clk_period;
Addr <= "0100010111011";
Trees_din <= "00000110000000000000000000000100";
wait for Clk_period;
Addr <= "0100010111100";
Trees_din <= "00000000000101100010010010101101";
wait for Clk_period;
Addr <= "0100010111101";
Trees_din <= "00000000000010110010010010101101";
wait for Clk_period;
Addr <= "0100010111110";
Trees_din <= "00000010000000000011111100010000";
wait for Clk_period;
Addr <= "0100010111111";
Trees_din <= "00000011000000000010000100001000";
wait for Clk_period;
Addr <= "0100011000000";
Trees_din <= "00000110000000000010010100000100";
wait for Clk_period;
Addr <= "0100011000001";
Trees_din <= "00000000001000100010010010101101";
wait for Clk_period;
Addr <= "0100011000010";
Trees_din <= "00000000000010100010010010101101";
wait for Clk_period;
Addr <= "0100011000011";
Trees_din <= "00000100000000000001100100000100";
wait for Clk_period;
Addr <= "0100011000100";
Trees_din <= "00000000000010100010010010101101";
wait for Clk_period;
Addr <= "0100011000101";
Trees_din <= "00000000001001000010010010101101";
wait for Clk_period;
Addr <= "0100011000110";
Trees_din <= "00000011000000000000111000001000";
wait for Clk_period;
Addr <= "0100011000111";
Trees_din <= "00000101000000000000100000000100";
wait for Clk_period;
Addr <= "0100011001000";
Trees_din <= "00000000010101000010010010101101";
wait for Clk_period;
Addr <= "0100011001001";
Trees_din <= "00000000010011000010010010101101";
wait for Clk_period;
Addr <= "0100011001010";
Trees_din <= "00000001000000000101111100000100";
wait for Clk_period;
Addr <= "0100011001011";
Trees_din <= "00000000010110110010010010101101";
wait for Clk_period;
Addr <= "0100011001100";
Trees_din <= "00000000010010000010010010101101";
wait for Clk_period;
Addr <= "0100011001101";
Trees_din <= "00000010000000000011100100100000";
wait for Clk_period;
Addr <= "0100011001110";
Trees_din <= "00000111000000000000011100010000";
wait for Clk_period;
Addr <= "0100011001111";
Trees_din <= "00000100000000000001011100001000";
wait for Clk_period;
Addr <= "0100011010000";
Trees_din <= "00000100000000000001010000000100";
wait for Clk_period;
Addr <= "0100011010001";
Trees_din <= "00000000000111110010010010101101";
wait for Clk_period;
Addr <= "0100011010010";
Trees_din <= "00000000000110010010010010101101";
wait for Clk_period;
Addr <= "0100011010011";
Trees_din <= "00000000000000000011100000000100";
wait for Clk_period;
Addr <= "0100011010100";
Trees_din <= "00000000010100110010010010101101";
wait for Clk_period;
Addr <= "0100011010101";
Trees_din <= "00000000000011110010010010101101";
wait for Clk_period;
Addr <= "0100011010110";
Trees_din <= "00000101000000000010110100001000";
wait for Clk_period;
Addr <= "0100011010111";
Trees_din <= "00000001000000000011100100000100";
wait for Clk_period;
Addr <= "0100011011000";
Trees_din <= "00000000000110000010010010101101";
wait for Clk_period;
Addr <= "0100011011001";
Trees_din <= "00000000000110000010010010101101";
wait for Clk_period;
Addr <= "0100011011010";
Trees_din <= "00000000000000000100010000000100";
wait for Clk_period;
Addr <= "0100011011011";
Trees_din <= "00000000011000110010010010101101";
wait for Clk_period;
Addr <= "0100011011100";
Trees_din <= "00000000010110000010010010101101";
wait for Clk_period;
Addr <= "0100011011101";
Trees_din <= "00000100000000000101110100010000";
wait for Clk_period;
Addr <= "0100011011110";
Trees_din <= "00000100000000000110001100001000";
wait for Clk_period;
Addr <= "0100011011111";
Trees_din <= "00000100000000000001110000000100";
wait for Clk_period;
Addr <= "0100011100000";
Trees_din <= "00000000011000000010010010101101";
wait for Clk_period;
Addr <= "0100011100001";
Trees_din <= "00000000011001000010010010101101";
wait for Clk_period;
Addr <= "0100011100010";
Trees_din <= "00000111000000000000110000000100";
wait for Clk_period;
Addr <= "0100011100011";
Trees_din <= "00000000000110010010010010101101";
wait for Clk_period;
Addr <= "0100011100100";
Trees_din <= "00000000001100110010010010101101";
wait for Clk_period;
Addr <= "0100011100101";
Trees_din <= "00000111000000000011101000001000";
wait for Clk_period;
Addr <= "0100011100110";
Trees_din <= "00000011000000000000111100000100";
wait for Clk_period;
Addr <= "0100011100111";
Trees_din <= "00000000001111000010010010101101";
wait for Clk_period;
Addr <= "0100011101000";
Trees_din <= "00000000010110000010010010101101";
wait for Clk_period;
Addr <= "0100011101001";
Trees_din <= "00000001000000000011011000000100";
wait for Clk_period;
Addr <= "0100011101010";
Trees_din <= "00000000010011100010010010101101";
wait for Clk_period;
Addr <= "0100011101011";
Trees_din <= "00000000001011110010010010101101";
wait for Clk_period;
Addr <= "0100011101100";
Trees_din <= "00000111000000000011010001000000";
wait for Clk_period;
Addr <= "0100011101101";
Trees_din <= "00000010000000000000010000100000";
wait for Clk_period;
Addr <= "0100011101110";
Trees_din <= "00000111000000000110010000010000";
wait for Clk_period;
Addr <= "0100011101111";
Trees_din <= "00000100000000000011111000001000";
wait for Clk_period;
Addr <= "0100011110000";
Trees_din <= "00000000000000000100001000000100";
wait for Clk_period;
Addr <= "0100011110001";
Trees_din <= "00000000010101110010010010101101";
wait for Clk_period;
Addr <= "0100011110010";
Trees_din <= "00000000010000010010010010101101";
wait for Clk_period;
Addr <= "0100011110011";
Trees_din <= "00000011000000000001100100000100";
wait for Clk_period;
Addr <= "0100011110100";
Trees_din <= "00000000000001000010010010101101";
wait for Clk_period;
Addr <= "0100011110101";
Trees_din <= "00000000001001010010010010101101";
wait for Clk_period;
Addr <= "0100011110110";
Trees_din <= "00000101000000000101111000001000";
wait for Clk_period;
Addr <= "0100011110111";
Trees_din <= "00000011000000000001110100000100";
wait for Clk_period;
Addr <= "0100011111000";
Trees_din <= "00000000001001110010010010101101";
wait for Clk_period;
Addr <= "0100011111001";
Trees_din <= "00000000000101110010010010101101";
wait for Clk_period;
Addr <= "0100011111010";
Trees_din <= "00000111000000000010101000000100";
wait for Clk_period;
Addr <= "0100011111011";
Trees_din <= "00000000010010000010010010101101";
wait for Clk_period;
Addr <= "0100011111100";
Trees_din <= "00000000001000000010010010101101";
wait for Clk_period;
Addr <= "0100011111101";
Trees_din <= "00000001000000000001100000010000";
wait for Clk_period;
Addr <= "0100011111110";
Trees_din <= "00000110000000000101111000001000";
wait for Clk_period;
Addr <= "0100011111111";
Trees_din <= "00000101000000000101110000000100";
wait for Clk_period;
Addr <= "0100100000000";
Trees_din <= "00000000000001000010010010101101";
wait for Clk_period;
Addr <= "0100100000001";
Trees_din <= "00000000001000100010010010101101";
wait for Clk_period;
Addr <= "0100100000010";
Trees_din <= "00000001000000000100110000000100";
wait for Clk_period;
Addr <= "0100100000011";
Trees_din <= "00000000001100110010010010101101";
wait for Clk_period;
Addr <= "0100100000100";
Trees_din <= "00000000000010000010010010101101";
wait for Clk_period;
Addr <= "0100100000101";
Trees_din <= "00000001000000000101110100001000";
wait for Clk_period;
Addr <= "0100100000110";
Trees_din <= "00000001000000000110001100000100";
wait for Clk_period;
Addr <= "0100100000111";
Trees_din <= "00000000010001100010010010101101";
wait for Clk_period;
Addr <= "0100100001000";
Trees_din <= "00000000000101010010010010101101";
wait for Clk_period;
Addr <= "0100100001001";
Trees_din <= "00000110000000000101011100000100";
wait for Clk_period;
Addr <= "0100100001010";
Trees_din <= "00000000010110000010010010101101";
wait for Clk_period;
Addr <= "0100100001011";
Trees_din <= "00000000000101110010010010101101";
wait for Clk_period;
Addr <= "0100100001100";
Trees_din <= "00000100000000000000101000100000";
wait for Clk_period;
Addr <= "0100100001101";
Trees_din <= "00000111000000000011101100010000";
wait for Clk_period;
Addr <= "0100100001110";
Trees_din <= "00000101000000000100010000001000";
wait for Clk_period;
Addr <= "0100100001111";
Trees_din <= "00000000000000000110001000000100";
wait for Clk_period;
Addr <= "0100100010000";
Trees_din <= "00000000000110110010010010101101";
wait for Clk_period;
Addr <= "0100100010001";
Trees_din <= "00000000010110100010010010101101";
wait for Clk_period;
Addr <= "0100100010010";
Trees_din <= "00000000000000000011100100000100";
wait for Clk_period;
Addr <= "0100100010011";
Trees_din <= "00000000001101110010010010101101";
wait for Clk_period;
Addr <= "0100100010100";
Trees_din <= "00000000010010000010010010101101";
wait for Clk_period;
Addr <= "0100100010101";
Trees_din <= "00000011000000000101001100001000";
wait for Clk_period;
Addr <= "0100100010110";
Trees_din <= "00000011000000000011100100000100";
wait for Clk_period;
Addr <= "0100100010111";
Trees_din <= "00000000010001110010010010101101";
wait for Clk_period;
Addr <= "0100100011000";
Trees_din <= "00000000000101100010010010101101";
wait for Clk_period;
Addr <= "0100100011001";
Trees_din <= "00000001000000000010100100000100";
wait for Clk_period;
Addr <= "0100100011010";
Trees_din <= "00000000010001100010010010101101";
wait for Clk_period;
Addr <= "0100100011011";
Trees_din <= "00000000010001100010010010101101";
wait for Clk_period;
Addr <= "0100100011100";
Trees_din <= "00000110000000000011000000010000";
wait for Clk_period;
Addr <= "0100100011101";
Trees_din <= "00000110000000000001101100001000";
wait for Clk_period;
Addr <= "0100100011110";
Trees_din <= "00000001000000000001101100000100";
wait for Clk_period;
Addr <= "0100100011111";
Trees_din <= "00000000001010000010010010101101";
wait for Clk_period;
Addr <= "0100100100000";
Trees_din <= "00000000000110010010010010101101";
wait for Clk_period;
Addr <= "0100100100001";
Trees_din <= "00000010000000000000100000000100";
wait for Clk_period;
Addr <= "0100100100010";
Trees_din <= "00000000010101110010010010101101";
wait for Clk_period;
Addr <= "0100100100011";
Trees_din <= "00000000001110100010010010101101";
wait for Clk_period;
Addr <= "0100100100100";
Trees_din <= "00000000000000000011101000001000";
wait for Clk_period;
Addr <= "0100100100101";
Trees_din <= "00000101000000000000111100000100";
wait for Clk_period;
Addr <= "0100100100110";
Trees_din <= "00000000010001010010010010101101";
wait for Clk_period;
Addr <= "0100100100111";
Trees_din <= "00000000000101110010010010101101";
wait for Clk_period;
Addr <= "0100100101000";
Trees_din <= "00000000000000000100101000000100";
wait for Clk_period;
Addr <= "0100100101001";
Trees_din <= "00000000001011100010010010101101";
wait for Clk_period;
Addr <= "0100100101010";
Trees_din <= "00000000001100110010010010101101";
wait for Clk_period;



----------tree 18-------------------

Addr <= "0100100101011";
Trees_din <= "00000001000000000011111110000000";
wait for Clk_period;
Addr <= "0100100101100";
Trees_din <= "00000100000000000001011001000000";
wait for Clk_period;
Addr <= "0100100101101";
Trees_din <= "00000000000000000100101000100000";
wait for Clk_period;
Addr <= "0100100101110";
Trees_din <= "00000110000000000010101000010000";
wait for Clk_period;
Addr <= "0100100101111";
Trees_din <= "00000101000000000000110000001000";
wait for Clk_period;
Addr <= "0100100110000";
Trees_din <= "00000010000000000010111100000100";
wait for Clk_period;
Addr <= "0100100110001";
Trees_din <= "00000000011000100010011010101001";
wait for Clk_period;
Addr <= "0100100110010";
Trees_din <= "00000000000111010010011010101001";
wait for Clk_period;
Addr <= "0100100110011";
Trees_din <= "00000100000000000000100100000100";
wait for Clk_period;
Addr <= "0100100110100";
Trees_din <= "00000000000101000010011010101001";
wait for Clk_period;
Addr <= "0100100110101";
Trees_din <= "00000000000011100010011010101001";
wait for Clk_period;
Addr <= "0100100110110";
Trees_din <= "00000000000000000010101000001000";
wait for Clk_period;
Addr <= "0100100110111";
Trees_din <= "00000111000000000010111100000100";
wait for Clk_period;
Addr <= "0100100111000";
Trees_din <= "00000000000000000010011010101001";
wait for Clk_period;
Addr <= "0100100111001";
Trees_din <= "00000000000101110010011010101001";
wait for Clk_period;
Addr <= "0100100111010";
Trees_din <= "00000100000000000011101100000100";
wait for Clk_period;
Addr <= "0100100111011";
Trees_din <= "00000000001110100010011010101001";
wait for Clk_period;
Addr <= "0100100111100";
Trees_din <= "00000000001010100010011010101001";
wait for Clk_period;
Addr <= "0100100111101";
Trees_din <= "00000011000000000001011100010000";
wait for Clk_period;
Addr <= "0100100111110";
Trees_din <= "00000101000000000000110000001000";
wait for Clk_period;
Addr <= "0100100111111";
Trees_din <= "00000010000000000101101100000100";
wait for Clk_period;
Addr <= "0100101000000";
Trees_din <= "00000000000011000010011010101001";
wait for Clk_period;
Addr <= "0100101000001";
Trees_din <= "00000000010111100010011010101001";
wait for Clk_period;
Addr <= "0100101000010";
Trees_din <= "00000000000000000000001100000100";
wait for Clk_period;
Addr <= "0100101000011";
Trees_din <= "00000000001100100010011010101001";
wait for Clk_period;
Addr <= "0100101000100";
Trees_din <= "00000000010101110010011010101001";
wait for Clk_period;
Addr <= "0100101000101";
Trees_din <= "00000110000000000100100000001000";
wait for Clk_period;
Addr <= "0100101000110";
Trees_din <= "00000010000000000000000000000100";
wait for Clk_period;
Addr <= "0100101000111";
Trees_din <= "00000000010010110010011010101001";
wait for Clk_period;
Addr <= "0100101001000";
Trees_din <= "00000000000011010010011010101001";
wait for Clk_period;
Addr <= "0100101001001";
Trees_din <= "00000111000000000000011000000100";
wait for Clk_period;
Addr <= "0100101001010";
Trees_din <= "00000000001010000010011010101001";
wait for Clk_period;
Addr <= "0100101001011";
Trees_din <= "00000000010101100010011010101001";
wait for Clk_period;
Addr <= "0100101001100";
Trees_din <= "00000101000000000000101100100000";
wait for Clk_period;
Addr <= "0100101001101";
Trees_din <= "00000100000000000001001000010000";
wait for Clk_period;
Addr <= "0100101001110";
Trees_din <= "00000010000000000000000100001000";
wait for Clk_period;
Addr <= "0100101001111";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "0100101010000";
Trees_din <= "00000000000001100010011010101001";
wait for Clk_period;
Addr <= "0100101010001";
Trees_din <= "00000000000000000010011010101001";
wait for Clk_period;
Addr <= "0100101010010";
Trees_din <= "00000100000000000001001100000100";
wait for Clk_period;
Addr <= "0100101010011";
Trees_din <= "00000000000101110010011010101001";
wait for Clk_period;
Addr <= "0100101010100";
Trees_din <= "00000000000011100010011010101001";
wait for Clk_period;
Addr <= "0100101010101";
Trees_din <= "00000001000000000000010000001000";
wait for Clk_period;
Addr <= "0100101010110";
Trees_din <= "00000001000000000001011000000100";
wait for Clk_period;
Addr <= "0100101010111";
Trees_din <= "00000000010011110010011010101001";
wait for Clk_period;
Addr <= "0100101011000";
Trees_din <= "00000000000001010010011010101001";
wait for Clk_period;
Addr <= "0100101011001";
Trees_din <= "00000000000000000100010000000100";
wait for Clk_period;
Addr <= "0100101011010";
Trees_din <= "00000000000101000010011010101001";
wait for Clk_period;
Addr <= "0100101011011";
Trees_din <= "00000000010011110010011010101001";
wait for Clk_period;
Addr <= "0100101011100";
Trees_din <= "00000101000000000100101000010000";
wait for Clk_period;
Addr <= "0100101011101";
Trees_din <= "00000101000000000100100100001000";
wait for Clk_period;
Addr <= "0100101011110";
Trees_din <= "00000110000000000100111000000100";
wait for Clk_period;
Addr <= "0100101011111";
Trees_din <= "00000000010101000010011010101001";
wait for Clk_period;
Addr <= "0100101100000";
Trees_din <= "00000000001000010010011010101001";
wait for Clk_period;
Addr <= "0100101100001";
Trees_din <= "00000000000000000000100000000100";
wait for Clk_period;
Addr <= "0100101100010";
Trees_din <= "00000000001111110010011010101001";
wait for Clk_period;
Addr <= "0100101100011";
Trees_din <= "00000000010110110010011010101001";
wait for Clk_period;
Addr <= "0100101100100";
Trees_din <= "00000100000000000010001000001000";
wait for Clk_period;
Addr <= "0100101100101";
Trees_din <= "00000011000000000001011000000100";
wait for Clk_period;
Addr <= "0100101100110";
Trees_din <= "00000000000101110010011010101001";
wait for Clk_period;
Addr <= "0100101100111";
Trees_din <= "00000000010101100010011010101001";
wait for Clk_period;
Addr <= "0100101101000";
Trees_din <= "00000001000000000101010100000100";
wait for Clk_period;
Addr <= "0100101101001";
Trees_din <= "00000000010100000010011010101001";
wait for Clk_period;
Addr <= "0100101101010";
Trees_din <= "00000000010000010010011010101001";
wait for Clk_period;
Addr <= "0100101101011";
Trees_din <= "00000010000000000100101001000000";
wait for Clk_period;
Addr <= "0100101101100";
Trees_din <= "00000010000000000010100100100000";
wait for Clk_period;
Addr <= "0100101101101";
Trees_din <= "00000101000000000110000000010000";
wait for Clk_period;
Addr <= "0100101101110";
Trees_din <= "00000111000000000011111000001000";
wait for Clk_period;
Addr <= "0100101101111";
Trees_din <= "00000010000000000001101100000100";
wait for Clk_period;
Addr <= "0100101110000";
Trees_din <= "00000000010000010010011010101001";
wait for Clk_period;
Addr <= "0100101110001";
Trees_din <= "00000000010000110010011010101001";
wait for Clk_period;
Addr <= "0100101110010";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0100101110011";
Trees_din <= "00000000000011000010011010101001";
wait for Clk_period;
Addr <= "0100101110100";
Trees_din <= "00000000000111100010011010101001";
wait for Clk_period;
Addr <= "0100101110101";
Trees_din <= "00000001000000000010110100001000";
wait for Clk_period;
Addr <= "0100101110110";
Trees_din <= "00000111000000000011000100000100";
wait for Clk_period;
Addr <= "0100101110111";
Trees_din <= "00000000000001010010011010101001";
wait for Clk_period;
Addr <= "0100101111000";
Trees_din <= "00000000001111000010011010101001";
wait for Clk_period;
Addr <= "0100101111001";
Trees_din <= "00000011000000000101001100000100";
wait for Clk_period;
Addr <= "0100101111010";
Trees_din <= "00000000000000010010011010101001";
wait for Clk_period;
Addr <= "0100101111011";
Trees_din <= "00000000010101100010011010101001";
wait for Clk_period;
Addr <= "0100101111100";
Trees_din <= "00000000000000000000110000010000";
wait for Clk_period;
Addr <= "0100101111101";
Trees_din <= "00000011000000000100011000001000";
wait for Clk_period;
Addr <= "0100101111110";
Trees_din <= "00000111000000000001011100000100";
wait for Clk_period;
Addr <= "0100101111111";
Trees_din <= "00000000010011010010011010101001";
wait for Clk_period;
Addr <= "0100110000000";
Trees_din <= "00000000000100110010011010101001";
wait for Clk_period;
Addr <= "0100110000001";
Trees_din <= "00000100000000000110010000000100";
wait for Clk_period;
Addr <= "0100110000010";
Trees_din <= "00000000010111100010011010101001";
wait for Clk_period;
Addr <= "0100110000011";
Trees_din <= "00000000000011010010011010101001";
wait for Clk_period;
Addr <= "0100110000100";
Trees_din <= "00000011000000000001001100001000";
wait for Clk_period;
Addr <= "0100110000101";
Trees_din <= "00000011000000000010100000000100";
wait for Clk_period;
Addr <= "0100110000110";
Trees_din <= "00000000000100110010011010101001";
wait for Clk_period;
Addr <= "0100110000111";
Trees_din <= "00000000000011000010011010101001";
wait for Clk_period;
Addr <= "0100110001000";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "0100110001001";
Trees_din <= "00000000001101110010011010101001";
wait for Clk_period;
Addr <= "0100110001010";
Trees_din <= "00000000001011010010011010101001";
wait for Clk_period;
Addr <= "0100110001011";
Trees_din <= "00000001000000000010000100100000";
wait for Clk_period;
Addr <= "0100110001100";
Trees_din <= "00000010000000000011110100010000";
wait for Clk_period;
Addr <= "0100110001101";
Trees_din <= "00000000000000000001100000001000";
wait for Clk_period;
Addr <= "0100110001110";
Trees_din <= "00000110000000000010011000000100";
wait for Clk_period;
Addr <= "0100110001111";
Trees_din <= "00000000010001100010011010101001";
wait for Clk_period;
Addr <= "0100110010000";
Trees_din <= "00000000001111010010011010101001";
wait for Clk_period;
Addr <= "0100110010001";
Trees_din <= "00000001000000000000111100000100";
wait for Clk_period;
Addr <= "0100110010010";
Trees_din <= "00000000001011110010011010101001";
wait for Clk_period;
Addr <= "0100110010011";
Trees_din <= "00000000010111100010011010101001";
wait for Clk_period;
Addr <= "0100110010100";
Trees_din <= "00000101000000000100100100001000";
wait for Clk_period;
Addr <= "0100110010101";
Trees_din <= "00000100000000000001001000000100";
wait for Clk_period;
Addr <= "0100110010110";
Trees_din <= "00000000001101100010011010101001";
wait for Clk_period;
Addr <= "0100110010111";
Trees_din <= "00000000010011010010011010101001";
wait for Clk_period;
Addr <= "0100110011000";
Trees_din <= "00000100000000000100001100000100";
wait for Clk_period;
Addr <= "0100110011001";
Trees_din <= "00000000000101010010011010101001";
wait for Clk_period;
Addr <= "0100110011010";
Trees_din <= "00000000010110000010011010101001";
wait for Clk_period;
Addr <= "0100110011011";
Trees_din <= "00000010000000000101010100010000";
wait for Clk_period;
Addr <= "0100110011100";
Trees_din <= "00000010000000000001000100001000";
wait for Clk_period;
Addr <= "0100110011101";
Trees_din <= "00000101000000000001101000000100";
wait for Clk_period;
Addr <= "0100110011110";
Trees_din <= "00000000011000100010011010101001";
wait for Clk_period;
Addr <= "0100110011111";
Trees_din <= "00000000000001100010011010101001";
wait for Clk_period;
Addr <= "0100110100000";
Trees_din <= "00000000000000000010000100000100";
wait for Clk_period;
Addr <= "0100110100001";
Trees_din <= "00000000000101000010011010101001";
wait for Clk_period;
Addr <= "0100110100010";
Trees_din <= "00000000001010000010011010101001";
wait for Clk_period;
Addr <= "0100110100011";
Trees_din <= "00000000000000000100000000001000";
wait for Clk_period;
Addr <= "0100110100100";
Trees_din <= "00000111000000000101011100000100";
wait for Clk_period;
Addr <= "0100110100101";
Trees_din <= "00000000000001110010011010101001";
wait for Clk_period;
Addr <= "0100110100110";
Trees_din <= "00000000010010000010011010101001";
wait for Clk_period;
Addr <= "0100110100111";
Trees_din <= "00000100000000000011000000000100";
wait for Clk_period;
Addr <= "0100110101000";
Trees_din <= "00000000010010110010011010101001";
wait for Clk_period;
Addr <= "0100110101001";
Trees_din <= "00000000010000110010011010101001";
wait for Clk_period;



----------tree 19-------------------

Addr <= "0100110101010";
Trees_din <= "00000101000000000000011010000000";
wait for Clk_period;
Addr <= "0100110101011";
Trees_din <= "00000110000000000100011101000000";
wait for Clk_period;
Addr <= "0100110101100";
Trees_din <= "00000100000000000011110000100000";
wait for Clk_period;
Addr <= "0100110101101";
Trees_din <= "00000011000000000010110000010000";
wait for Clk_period;
Addr <= "0100110101110";
Trees_din <= "00000101000000000011110100001000";
wait for Clk_period;
Addr <= "0100110101111";
Trees_din <= "00000011000000000011001100000100";
wait for Clk_period;
Addr <= "0100110110000";
Trees_din <= "00000000010010110010100010100101";
wait for Clk_period;
Addr <= "0100110110001";
Trees_din <= "00000000001100100010100010100101";
wait for Clk_period;
Addr <= "0100110110010";
Trees_din <= "00000011000000000010100100000100";
wait for Clk_period;
Addr <= "0100110110011";
Trees_din <= "00000000001001100010100010100101";
wait for Clk_period;
Addr <= "0100110110100";
Trees_din <= "00000000010011110010100010100101";
wait for Clk_period;
Addr <= "0100110110101";
Trees_din <= "00000000000000000001000100001000";
wait for Clk_period;
Addr <= "0100110110110";
Trees_din <= "00000110000000000101100100000100";
wait for Clk_period;
Addr <= "0100110110111";
Trees_din <= "00000000010001000010100010100101";
wait for Clk_period;
Addr <= "0100110111000";
Trees_din <= "00000000000110110010100010100101";
wait for Clk_period;
Addr <= "0100110111001";
Trees_din <= "00000010000000000010111000000100";
wait for Clk_period;
Addr <= "0100110111010";
Trees_din <= "00000000000011100010100010100101";
wait for Clk_period;
Addr <= "0100110111011";
Trees_din <= "00000000000101010010100010100101";
wait for Clk_period;
Addr <= "0100110111100";
Trees_din <= "00000000000000000110000100010000";
wait for Clk_period;
Addr <= "0100110111101";
Trees_din <= "00000110000000000001000100001000";
wait for Clk_period;
Addr <= "0100110111110";
Trees_din <= "00000101000000000011011000000100";
wait for Clk_period;
Addr <= "0100110111111";
Trees_din <= "00000000001011100010100010100101";
wait for Clk_period;
Addr <= "0100111000000";
Trees_din <= "00000000000101010010100010100101";
wait for Clk_period;
Addr <= "0100111000001";
Trees_din <= "00000011000000000001110100000100";
wait for Clk_period;
Addr <= "0100111000010";
Trees_din <= "00000000000011010010100010100101";
wait for Clk_period;
Addr <= "0100111000011";
Trees_din <= "00000000001001010010100010100101";
wait for Clk_period;
Addr <= "0100111000100";
Trees_din <= "00000001000000000110001100001000";
wait for Clk_period;
Addr <= "0100111000101";
Trees_din <= "00000100000000000001100100000100";
wait for Clk_period;
Addr <= "0100111000110";
Trees_din <= "00000000001010010010100010100101";
wait for Clk_period;
Addr <= "0100111000111";
Trees_din <= "00000000001010100010100010100101";
wait for Clk_period;
Addr <= "0100111001000";
Trees_din <= "00000110000000000101100000000100";
wait for Clk_period;
Addr <= "0100111001001";
Trees_din <= "00000000010111010010100010100101";
wait for Clk_period;
Addr <= "0100111001010";
Trees_din <= "00000000000000100010100010100101";
wait for Clk_period;
Addr <= "0100111001011";
Trees_din <= "00000111000000000011011000100000";
wait for Clk_period;
Addr <= "0100111001100";
Trees_din <= "00000000000000000100111100010000";
wait for Clk_period;
Addr <= "0100111001101";
Trees_din <= "00000000000000000000010100001000";
wait for Clk_period;
Addr <= "0100111001110";
Trees_din <= "00000111000000000010100100000100";
wait for Clk_period;
Addr <= "0100111001111";
Trees_din <= "00000000010110010010100010100101";
wait for Clk_period;
Addr <= "0100111010000";
Trees_din <= "00000000000111000010100010100101";
wait for Clk_period;
Addr <= "0100111010001";
Trees_din <= "00000011000000000001000100000100";
wait for Clk_period;
Addr <= "0100111010010";
Trees_din <= "00000000010110110010100010100101";
wait for Clk_period;
Addr <= "0100111010011";
Trees_din <= "00000000010110110010100010100101";
wait for Clk_period;
Addr <= "0100111010100";
Trees_din <= "00000100000000000011011000001000";
wait for Clk_period;
Addr <= "0100111010101";
Trees_din <= "00000001000000000011001000000100";
wait for Clk_period;
Addr <= "0100111010110";
Trees_din <= "00000000001001110010100010100101";
wait for Clk_period;
Addr <= "0100111010111";
Trees_din <= "00000000000000110010100010100101";
wait for Clk_period;
Addr <= "0100111011000";
Trees_din <= "00000100000000000010100100000100";
wait for Clk_period;
Addr <= "0100111011001";
Trees_din <= "00000000010010100010100010100101";
wait for Clk_period;
Addr <= "0100111011010";
Trees_din <= "00000000000111010010100010100101";
wait for Clk_period;
Addr <= "0100111011011";
Trees_din <= "00000100000000000011000100010000";
wait for Clk_period;
Addr <= "0100111011100";
Trees_din <= "00000010000000000001111000001000";
wait for Clk_period;
Addr <= "0100111011101";
Trees_din <= "00000100000000000001011100000100";
wait for Clk_period;
Addr <= "0100111011110";
Trees_din <= "00000000010001100010100010100101";
wait for Clk_period;
Addr <= "0100111011111";
Trees_din <= "00000000001010100010100010100101";
wait for Clk_period;
Addr <= "0100111100000";
Trees_din <= "00000101000000000101110000000100";
wait for Clk_period;
Addr <= "0100111100001";
Trees_din <= "00000000000111000010100010100101";
wait for Clk_period;
Addr <= "0100111100010";
Trees_din <= "00000000001000010010100010100101";
wait for Clk_period;
Addr <= "0100111100011";
Trees_din <= "00000001000000000001100100001000";
wait for Clk_period;
Addr <= "0100111100100";
Trees_din <= "00000000000000000010110100000100";
wait for Clk_period;
Addr <= "0100111100101";
Trees_din <= "00000000001101110010100010100101";
wait for Clk_period;
Addr <= "0100111100110";
Trees_din <= "00000000000100100010100010100101";
wait for Clk_period;
Addr <= "0100111100111";
Trees_din <= "00000100000000000000011000000100";
wait for Clk_period;
Addr <= "0100111101000";
Trees_din <= "00000000001011010010100010100101";
wait for Clk_period;
Addr <= "0100111101001";
Trees_din <= "00000000010100010010100010100101";
wait for Clk_period;
Addr <= "0100111101010";
Trees_din <= "00000111000000000001001101000000";
wait for Clk_period;
Addr <= "0100111101011";
Trees_din <= "00000001000000000100001000100000";
wait for Clk_period;
Addr <= "0100111101100";
Trees_din <= "00000110000000000011100000010000";
wait for Clk_period;
Addr <= "0100111101101";
Trees_din <= "00000000000000000000000000001000";
wait for Clk_period;
Addr <= "0100111101110";
Trees_din <= "00000000000000000100101100000100";
wait for Clk_period;
Addr <= "0100111101111";
Trees_din <= "00000000000111010010100010100101";
wait for Clk_period;
Addr <= "0100111110000";
Trees_din <= "00000000010101000010100010100101";
wait for Clk_period;
Addr <= "0100111110001";
Trees_din <= "00000111000000000011101000000100";
wait for Clk_period;
Addr <= "0100111110010";
Trees_din <= "00000000010011110010100010100101";
wait for Clk_period;
Addr <= "0100111110011";
Trees_din <= "00000000000100010010100010100101";
wait for Clk_period;
Addr <= "0100111110100";
Trees_din <= "00000010000000000001000100001000";
wait for Clk_period;
Addr <= "0100111110101";
Trees_din <= "00000110000000000100101100000100";
wait for Clk_period;
Addr <= "0100111110110";
Trees_din <= "00000000001010010010100010100101";
wait for Clk_period;
Addr <= "0100111110111";
Trees_din <= "00000000001110100010100010100101";
wait for Clk_period;
Addr <= "0100111111000";
Trees_din <= "00000001000000000010011100000100";
wait for Clk_period;
Addr <= "0100111111001";
Trees_din <= "00000000010100110010100010100101";
wait for Clk_period;
Addr <= "0100111111010";
Trees_din <= "00000000001111000010100010100101";
wait for Clk_period;
Addr <= "0100111111011";
Trees_din <= "00000100000000000010000000010000";
wait for Clk_period;
Addr <= "0100111111100";
Trees_din <= "00000001000000000110000100001000";
wait for Clk_period;
Addr <= "0100111111101";
Trees_din <= "00000101000000000101111100000100";
wait for Clk_period;
Addr <= "0100111111110";
Trees_din <= "00000000001111010010100010100101";
wait for Clk_period;
Addr <= "0100111111111";
Trees_din <= "00000000000000110010100010100101";
wait for Clk_period;
Addr <= "0101000000000";
Trees_din <= "00000010000000000101111000000100";
wait for Clk_period;
Addr <= "0101000000001";
Trees_din <= "00000000000011010010100010100101";
wait for Clk_period;
Addr <= "0101000000010";
Trees_din <= "00000000000110000010100010100101";
wait for Clk_period;
Addr <= "0101000000011";
Trees_din <= "00000000000000000010011000001000";
wait for Clk_period;
Addr <= "0101000000100";
Trees_din <= "00000101000000000001110100000100";
wait for Clk_period;
Addr <= "0101000000101";
Trees_din <= "00000000000111010010100010100101";
wait for Clk_period;
Addr <= "0101000000110";
Trees_din <= "00000000010010000010100010100101";
wait for Clk_period;
Addr <= "0101000000111";
Trees_din <= "00000101000000000011000100000100";
wait for Clk_period;
Addr <= "0101000001000";
Trees_din <= "00000000000111110010100010100101";
wait for Clk_period;
Addr <= "0101000001001";
Trees_din <= "00000000001000100010100010100101";
wait for Clk_period;
Addr <= "0101000001010";
Trees_din <= "00000110000000000001011100100000";
wait for Clk_period;
Addr <= "0101000001011";
Trees_din <= "00000110000000000010100000010000";
wait for Clk_period;
Addr <= "0101000001100";
Trees_din <= "00000011000000000000111000001000";
wait for Clk_period;
Addr <= "0101000001101";
Trees_din <= "00000001000000000100010100000100";
wait for Clk_period;
Addr <= "0101000001110";
Trees_din <= "00000000000000100010100010100101";
wait for Clk_period;
Addr <= "0101000001111";
Trees_din <= "00000000000011110010100010100101";
wait for Clk_period;
Addr <= "0101000010000";
Trees_din <= "00000100000000000011101100000100";
wait for Clk_period;
Addr <= "0101000010001";
Trees_din <= "00000000001011100010100010100101";
wait for Clk_period;
Addr <= "0101000010010";
Trees_din <= "00000000000111100010100010100101";
wait for Clk_period;
Addr <= "0101000010011";
Trees_din <= "00000101000000000001001100001000";
wait for Clk_period;
Addr <= "0101000010100";
Trees_din <= "00000110000000000010000100000100";
wait for Clk_period;
Addr <= "0101000010101";
Trees_din <= "00000000010000000010100010100101";
wait for Clk_period;
Addr <= "0101000010110";
Trees_din <= "00000000000001110010100010100101";
wait for Clk_period;
Addr <= "0101000010111";
Trees_din <= "00000100000000000000010000000100";
wait for Clk_period;
Addr <= "0101000011000";
Trees_din <= "00000000001000010010100010100101";
wait for Clk_period;
Addr <= "0101000011001";
Trees_din <= "00000000010011110010100010100101";
wait for Clk_period;
Addr <= "0101000011010";
Trees_din <= "00000100000000000001010100010000";
wait for Clk_period;
Addr <= "0101000011011";
Trees_din <= "00000101000000000011000100001000";
wait for Clk_period;
Addr <= "0101000011100";
Trees_din <= "00000000000000000010110000000100";
wait for Clk_period;
Addr <= "0101000011101";
Trees_din <= "00000000010011100010100010100101";
wait for Clk_period;
Addr <= "0101000011110";
Trees_din <= "00000000000011100010100010100101";
wait for Clk_period;
Addr <= "0101000011111";
Trees_din <= "00000101000000000101101100000100";
wait for Clk_period;
Addr <= "0101000100000";
Trees_din <= "00000000000011110010100010100101";
wait for Clk_period;
Addr <= "0101000100001";
Trees_din <= "00000000001101100010100010100101";
wait for Clk_period;
Addr <= "0101000100010";
Trees_din <= "00000100000000000000011000001000";
wait for Clk_period;
Addr <= "0101000100011";
Trees_din <= "00000000000000000010001100000100";
wait for Clk_period;
Addr <= "0101000100100";
Trees_din <= "00000000010101010010100010100101";
wait for Clk_period;
Addr <= "0101000100101";
Trees_din <= "00000000010110100010100010100101";
wait for Clk_period;
Addr <= "0101000100110";
Trees_din <= "00000011000000000010101000000100";
wait for Clk_period;
Addr <= "0101000100111";
Trees_din <= "00000000001110010010100010100101";
wait for Clk_period;
Addr <= "0101000101000";
Trees_din <= "00000000001111010010100010100101";
wait for Clk_period;



----------tree 20-------------------

Addr <= "0101000101001";
Trees_din <= "00000110000000000001101110000000";
wait for Clk_period;
Addr <= "0101000101010";
Trees_din <= "00000100000000000101101101000000";
wait for Clk_period;
Addr <= "0101000101011";
Trees_din <= "00000011000000000001001000100000";
wait for Clk_period;
Addr <= "0101000101100";
Trees_din <= "00000011000000000100010100010000";
wait for Clk_period;
Addr <= "0101000101101";
Trees_din <= "00000000000000000000111100001000";
wait for Clk_period;
Addr <= "0101000101110";
Trees_din <= "00000111000000000000011000000100";
wait for Clk_period;
Addr <= "0101000101111";
Trees_din <= "00000000000001100010101010100001";
wait for Clk_period;
Addr <= "0101000110000";
Trees_din <= "00000000010110100010101010100001";
wait for Clk_period;
Addr <= "0101000110001";
Trees_din <= "00000010000000000101001000000100";
wait for Clk_period;
Addr <= "0101000110010";
Trees_din <= "00000000010100010010101010100001";
wait for Clk_period;
Addr <= "0101000110011";
Trees_din <= "00000000000001010010101010100001";
wait for Clk_period;
Addr <= "0101000110100";
Trees_din <= "00000000000000000100100100001000";
wait for Clk_period;
Addr <= "0101000110101";
Trees_din <= "00000011000000000000110000000100";
wait for Clk_period;
Addr <= "0101000110110";
Trees_din <= "00000000010010010010101010100001";
wait for Clk_period;
Addr <= "0101000110111";
Trees_din <= "00000000001110000010101010100001";
wait for Clk_period;
Addr <= "0101000111000";
Trees_din <= "00000011000000000010001100000100";
wait for Clk_period;
Addr <= "0101000111001";
Trees_din <= "00000000001000110010101010100001";
wait for Clk_period;
Addr <= "0101000111010";
Trees_din <= "00000000010000010010101010100001";
wait for Clk_period;
Addr <= "0101000111011";
Trees_din <= "00000101000000000011100100010000";
wait for Clk_period;
Addr <= "0101000111100";
Trees_din <= "00000110000000000001011100001000";
wait for Clk_period;
Addr <= "0101000111101";
Trees_din <= "00000010000000000000000000000100";
wait for Clk_period;
Addr <= "0101000111110";
Trees_din <= "00000000000100100010101010100001";
wait for Clk_period;
Addr <= "0101000111111";
Trees_din <= "00000000010010010010101010100001";
wait for Clk_period;
Addr <= "0101001000000";
Trees_din <= "00000000000000000010001100000100";
wait for Clk_period;
Addr <= "0101001000001";
Trees_din <= "00000000001011000010101010100001";
wait for Clk_period;
Addr <= "0101001000010";
Trees_din <= "00000000000110110010101010100001";
wait for Clk_period;
Addr <= "0101001000011";
Trees_din <= "00000110000000000010110100001000";
wait for Clk_period;
Addr <= "0101001000100";
Trees_din <= "00000001000000000110001100000100";
wait for Clk_period;
Addr <= "0101001000101";
Trees_din <= "00000000000000010010101010100001";
wait for Clk_period;
Addr <= "0101001000110";
Trees_din <= "00000000001110100010101010100001";
wait for Clk_period;
Addr <= "0101001000111";
Trees_din <= "00000101000000000001100100000100";
wait for Clk_period;
Addr <= "0101001001000";
Trees_din <= "00000000011001000010101010100001";
wait for Clk_period;
Addr <= "0101001001001";
Trees_din <= "00000000000110010010101010100001";
wait for Clk_period;
Addr <= "0101001001010";
Trees_din <= "00000000000000000010001000100000";
wait for Clk_period;
Addr <= "0101001001011";
Trees_din <= "00000111000000000011111000010000";
wait for Clk_period;
Addr <= "0101001001100";
Trees_din <= "00000101000000000001110000001000";
wait for Clk_period;
Addr <= "0101001001101";
Trees_din <= "00000111000000000001111100000100";
wait for Clk_period;
Addr <= "0101001001110";
Trees_din <= "00000000000100100010101010100001";
wait for Clk_period;
Addr <= "0101001001111";
Trees_din <= "00000000010000100010101010100001";
wait for Clk_period;
Addr <= "0101001010000";
Trees_din <= "00000110000000000010000000000100";
wait for Clk_period;
Addr <= "0101001010001";
Trees_din <= "00000000010001010010101010100001";
wait for Clk_period;
Addr <= "0101001010010";
Trees_din <= "00000000001010110010101010100001";
wait for Clk_period;
Addr <= "0101001010011";
Trees_din <= "00000000000000000100011000001000";
wait for Clk_period;
Addr <= "0101001010100";
Trees_din <= "00000001000000000011100000000100";
wait for Clk_period;
Addr <= "0101001010101";
Trees_din <= "00000000010001110010101010100001";
wait for Clk_period;
Addr <= "0101001010110";
Trees_din <= "00000000000010100010101010100001";
wait for Clk_period;
Addr <= "0101001010111";
Trees_din <= "00000010000000000101010100000100";
wait for Clk_period;
Addr <= "0101001011000";
Trees_din <= "00000000000011100010101010100001";
wait for Clk_period;
Addr <= "0101001011001";
Trees_din <= "00000000001000100010101010100001";
wait for Clk_period;
Addr <= "0101001011010";
Trees_din <= "00000111000000000110001000010000";
wait for Clk_period;
Addr <= "0101001011011";
Trees_din <= "00000100000000000001000100001000";
wait for Clk_period;
Addr <= "0101001011100";
Trees_din <= "00000111000000000100100000000100";
wait for Clk_period;
Addr <= "0101001011101";
Trees_din <= "00000000000000000010101010100001";
wait for Clk_period;
Addr <= "0101001011110";
Trees_din <= "00000000001101000010101010100001";
wait for Clk_period;
Addr <= "0101001011111";
Trees_din <= "00000011000000000000100000000100";
wait for Clk_period;
Addr <= "0101001100000";
Trees_din <= "00000000010110010010101010100001";
wait for Clk_period;
Addr <= "0101001100001";
Trees_din <= "00000000000100000010101010100001";
wait for Clk_period;
Addr <= "0101001100010";
Trees_din <= "00000101000000000001000100001000";
wait for Clk_period;
Addr <= "0101001100011";
Trees_din <= "00000101000000000010011100000100";
wait for Clk_period;
Addr <= "0101001100100";
Trees_din <= "00000000000011100010101010100001";
wait for Clk_period;
Addr <= "0101001100101";
Trees_din <= "00000000001111110010101010100001";
wait for Clk_period;
Addr <= "0101001100110";
Trees_din <= "00000010000000000101110000000100";
wait for Clk_period;
Addr <= "0101001100111";
Trees_din <= "00000000001010000010101010100001";
wait for Clk_period;
Addr <= "0101001101000";
Trees_din <= "00000000000100010010101010100001";
wait for Clk_period;
Addr <= "0101001101001";
Trees_din <= "00000101000000000001100001000000";
wait for Clk_period;
Addr <= "0101001101010";
Trees_din <= "00000110000000000000100000100000";
wait for Clk_period;
Addr <= "0101001101011";
Trees_din <= "00000001000000000110000100010000";
wait for Clk_period;
Addr <= "0101001101100";
Trees_din <= "00000101000000000000110100001000";
wait for Clk_period;
Addr <= "0101001101101";
Trees_din <= "00000000000000000100111000000100";
wait for Clk_period;
Addr <= "0101001101110";
Trees_din <= "00000000010011010010101010100001";
wait for Clk_period;
Addr <= "0101001101111";
Trees_din <= "00000000010111110010101010100001";
wait for Clk_period;
Addr <= "0101001110000";
Trees_din <= "00000101000000000010011000000100";
wait for Clk_period;
Addr <= "0101001110001";
Trees_din <= "00000000010110010010101010100001";
wait for Clk_period;
Addr <= "0101001110010";
Trees_din <= "00000000001000110010101010100001";
wait for Clk_period;
Addr <= "0101001110011";
Trees_din <= "00000010000000000011111000001000";
wait for Clk_period;
Addr <= "0101001110100";
Trees_din <= "00000000000000000011100000000100";
wait for Clk_period;
Addr <= "0101001110101";
Trees_din <= "00000000011001000010101010100001";
wait for Clk_period;
Addr <= "0101001110110";
Trees_din <= "00000000000000000010101010100001";
wait for Clk_period;
Addr <= "0101001110111";
Trees_din <= "00000100000000000000010000000100";
wait for Clk_period;
Addr <= "0101001111000";
Trees_din <= "00000000001010000010101010100001";
wait for Clk_period;
Addr <= "0101001111001";
Trees_din <= "00000000000011110010101010100001";
wait for Clk_period;
Addr <= "0101001111010";
Trees_din <= "00000010000000000000011000010000";
wait for Clk_period;
Addr <= "0101001111011";
Trees_din <= "00000110000000000000010100001000";
wait for Clk_period;
Addr <= "0101001111100";
Trees_din <= "00000101000000000000010100000100";
wait for Clk_period;
Addr <= "0101001111101";
Trees_din <= "00000000000111110010101010100001";
wait for Clk_period;
Addr <= "0101001111110";
Trees_din <= "00000000000010100010101010100001";
wait for Clk_period;
Addr <= "0101001111111";
Trees_din <= "00000100000000000101011000000100";
wait for Clk_period;
Addr <= "0101010000000";
Trees_din <= "00000000000010110010101010100001";
wait for Clk_period;
Addr <= "0101010000001";
Trees_din <= "00000000010000100010101010100001";
wait for Clk_period;
Addr <= "0101010000010";
Trees_din <= "00000110000000000001000000001000";
wait for Clk_period;
Addr <= "0101010000011";
Trees_din <= "00000111000000000000011000000100";
wait for Clk_period;
Addr <= "0101010000100";
Trees_din <= "00000000000010000010101010100001";
wait for Clk_period;
Addr <= "0101010000101";
Trees_din <= "00000000000111100010101010100001";
wait for Clk_period;
Addr <= "0101010000110";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "0101010000111";
Trees_din <= "00000000010101000010101010100001";
wait for Clk_period;
Addr <= "0101010001000";
Trees_din <= "00000000000110010010101010100001";
wait for Clk_period;
Addr <= "0101010001001";
Trees_din <= "00000100000000000101100000100000";
wait for Clk_period;
Addr <= "0101010001010";
Trees_din <= "00000111000000000100010000010000";
wait for Clk_period;
Addr <= "0101010001011";
Trees_din <= "00000010000000000011011100001000";
wait for Clk_period;
Addr <= "0101010001100";
Trees_din <= "00000010000000000000110100000100";
wait for Clk_period;
Addr <= "0101010001101";
Trees_din <= "00000000011000010010101010100001";
wait for Clk_period;
Addr <= "0101010001110";
Trees_din <= "00000000001011100010101010100001";
wait for Clk_period;
Addr <= "0101010001111";
Trees_din <= "00000101000000000000010000000100";
wait for Clk_period;
Addr <= "0101010010000";
Trees_din <= "00000000001011100010101010100001";
wait for Clk_period;
Addr <= "0101010010001";
Trees_din <= "00000000010111010010101010100001";
wait for Clk_period;
Addr <= "0101010010010";
Trees_din <= "00000000000000000011000000001000";
wait for Clk_period;
Addr <= "0101010010011";
Trees_din <= "00000111000000000101110100000100";
wait for Clk_period;
Addr <= "0101010010100";
Trees_din <= "00000000001100110010101010100001";
wait for Clk_period;
Addr <= "0101010010101";
Trees_din <= "00000000001001100010101010100001";
wait for Clk_period;
Addr <= "0101010010110";
Trees_din <= "00000111000000000011111100000100";
wait for Clk_period;
Addr <= "0101010010111";
Trees_din <= "00000000001111100010101010100001";
wait for Clk_period;
Addr <= "0101010011000";
Trees_din <= "00000000000101000010101010100001";
wait for Clk_period;
Addr <= "0101010011001";
Trees_din <= "00000100000000000010101100010000";
wait for Clk_period;
Addr <= "0101010011010";
Trees_din <= "00000000000000000011011100001000";
wait for Clk_period;
Addr <= "0101010011011";
Trees_din <= "00000111000000000000000000000100";
wait for Clk_period;
Addr <= "0101010011100";
Trees_din <= "00000000000111110010101010100001";
wait for Clk_period;
Addr <= "0101010011101";
Trees_din <= "00000000000101000010101010100001";
wait for Clk_period;
Addr <= "0101010011110";
Trees_din <= "00000010000000000110001000000100";
wait for Clk_period;
Addr <= "0101010011111";
Trees_din <= "00000000000101010010101010100001";
wait for Clk_period;
Addr <= "0101010100000";
Trees_din <= "00000000011000110010101010100001";
wait for Clk_period;
Addr <= "0101010100001";
Trees_din <= "00000100000000000010001100001000";
wait for Clk_period;
Addr <= "0101010100010";
Trees_din <= "00000111000000000100100100000100";
wait for Clk_period;
Addr <= "0101010100011";
Trees_din <= "00000000001011110010101010100001";
wait for Clk_period;
Addr <= "0101010100100";
Trees_din <= "00000000010110100010101010100001";
wait for Clk_period;
Addr <= "0101010100101";
Trees_din <= "00000010000000000001111100000100";
wait for Clk_period;
Addr <= "0101010100110";
Trees_din <= "00000000011000110010101010100001";
wait for Clk_period;
Addr <= "0101010100111";
Trees_din <= "00000000011000010010101010100001";
wait for Clk_period;



----------tree 21-------------------

Addr <= "0101010101000";
Trees_din <= "00000110000000000011001110000000";
wait for Clk_period;
Addr <= "0101010101001";
Trees_din <= "00000000000000000001000101000000";
wait for Clk_period;
Addr <= "0101010101010";
Trees_din <= "00000110000000000100110000100000";
wait for Clk_period;
Addr <= "0101010101011";
Trees_din <= "00000011000000000000011100010000";
wait for Clk_period;
Addr <= "0101010101100";
Trees_din <= "00000101000000000011010100001000";
wait for Clk_period;
Addr <= "0101010101101";
Trees_din <= "00000001000000000000111100000100";
wait for Clk_period;
Addr <= "0101010101110";
Trees_din <= "00000000001100010010110010011101";
wait for Clk_period;
Addr <= "0101010101111";
Trees_din <= "00000000001101110010110010011101";
wait for Clk_period;
Addr <= "0101010110000";
Trees_din <= "00000011000000000011101100000100";
wait for Clk_period;
Addr <= "0101010110001";
Trees_din <= "00000000000011010010110010011101";
wait for Clk_period;
Addr <= "0101010110010";
Trees_din <= "00000000000011110010110010011101";
wait for Clk_period;
Addr <= "0101010110011";
Trees_din <= "00000101000000000101010000001000";
wait for Clk_period;
Addr <= "0101010110100";
Trees_din <= "00000111000000000101100000000100";
wait for Clk_period;
Addr <= "0101010110101";
Trees_din <= "00000000011001000010110010011101";
wait for Clk_period;
Addr <= "0101010110110";
Trees_din <= "00000000001110100010110010011101";
wait for Clk_period;
Addr <= "0101010110111";
Trees_din <= "00000001000000000010011000000100";
wait for Clk_period;
Addr <= "0101010111000";
Trees_din <= "00000000001100100010110010011101";
wait for Clk_period;
Addr <= "0101010111001";
Trees_din <= "00000000001100110010110010011101";
wait for Clk_period;
Addr <= "0101010111010";
Trees_din <= "00000101000000000011000100010000";
wait for Clk_period;
Addr <= "0101010111011";
Trees_din <= "00000101000000000011100000001000";
wait for Clk_period;
Addr <= "0101010111100";
Trees_din <= "00000101000000000001100000000100";
wait for Clk_period;
Addr <= "0101010111101";
Trees_din <= "00000000000011000010110010011101";
wait for Clk_period;
Addr <= "0101010111110";
Trees_din <= "00000000000001000010110010011101";
wait for Clk_period;
Addr <= "0101010111111";
Trees_din <= "00000001000000000011001000000100";
wait for Clk_period;
Addr <= "0101011000000";
Trees_din <= "00000000000001100010110010011101";
wait for Clk_period;
Addr <= "0101011000001";
Trees_din <= "00000000011000100010110010011101";
wait for Clk_period;
Addr <= "0101011000010";
Trees_din <= "00000000000000000101100100001000";
wait for Clk_period;
Addr <= "0101011000011";
Trees_din <= "00000010000000000010001000000100";
wait for Clk_period;
Addr <= "0101011000100";
Trees_din <= "00000000001101110010110010011101";
wait for Clk_period;
Addr <= "0101011000101";
Trees_din <= "00000000000011100010110010011101";
wait for Clk_period;
Addr <= "0101011000110";
Trees_din <= "00000100000000000100011000000100";
wait for Clk_period;
Addr <= "0101011000111";
Trees_din <= "00000000000101010010110010011101";
wait for Clk_period;
Addr <= "0101011001000";
Trees_din <= "00000000010011010010110010011101";
wait for Clk_period;
Addr <= "0101011001001";
Trees_din <= "00000101000000000001110000100000";
wait for Clk_period;
Addr <= "0101011001010";
Trees_din <= "00000100000000000000110100010000";
wait for Clk_period;
Addr <= "0101011001011";
Trees_din <= "00000101000000000001000000001000";
wait for Clk_period;
Addr <= "0101011001100";
Trees_din <= "00000111000000000010101000000100";
wait for Clk_period;
Addr <= "0101011001101";
Trees_din <= "00000000010110010010110010011101";
wait for Clk_period;
Addr <= "0101011001110";
Trees_din <= "00000000001101010010110010011101";
wait for Clk_period;
Addr <= "0101011001111";
Trees_din <= "00000000000000000000100000000100";
wait for Clk_period;
Addr <= "0101011010000";
Trees_din <= "00000000001111100010110010011101";
wait for Clk_period;
Addr <= "0101011010001";
Trees_din <= "00000000000100110010110010011101";
wait for Clk_period;
Addr <= "0101011010010";
Trees_din <= "00000110000000000011101100001000";
wait for Clk_period;
Addr <= "0101011010011";
Trees_din <= "00000100000000000110000000000100";
wait for Clk_period;
Addr <= "0101011010100";
Trees_din <= "00000000010111100010110010011101";
wait for Clk_period;
Addr <= "0101011010101";
Trees_din <= "00000000010100110010110010011101";
wait for Clk_period;
Addr <= "0101011010110";
Trees_din <= "00000100000000000001011000000100";
wait for Clk_period;
Addr <= "0101011010111";
Trees_din <= "00000000000000100010110010011101";
wait for Clk_period;
Addr <= "0101011011000";
Trees_din <= "00000000010010000010110010011101";
wait for Clk_period;
Addr <= "0101011011001";
Trees_din <= "00000111000000000001100000010000";
wait for Clk_period;
Addr <= "0101011011010";
Trees_din <= "00000000000000000100101000001000";
wait for Clk_period;
Addr <= "0101011011011";
Trees_din <= "00000111000000000010010000000100";
wait for Clk_period;
Addr <= "0101011011100";
Trees_din <= "00000000000010000010110010011101";
wait for Clk_period;
Addr <= "0101011011101";
Trees_din <= "00000000010000110010110010011101";
wait for Clk_period;
Addr <= "0101011011110";
Trees_din <= "00000000000000000010110000000100";
wait for Clk_period;
Addr <= "0101011011111";
Trees_din <= "00000000000100100010110010011101";
wait for Clk_period;
Addr <= "0101011100000";
Trees_din <= "00000000000001100010110010011101";
wait for Clk_period;
Addr <= "0101011100001";
Trees_din <= "00000001000000000000011000001000";
wait for Clk_period;
Addr <= "0101011100010";
Trees_din <= "00000101000000000011110000000100";
wait for Clk_period;
Addr <= "0101011100011";
Trees_din <= "00000000010110100010110010011101";
wait for Clk_period;
Addr <= "0101011100100";
Trees_din <= "00000000000011010010110010011101";
wait for Clk_period;
Addr <= "0101011100101";
Trees_din <= "00000001000000000100001000000100";
wait for Clk_period;
Addr <= "0101011100110";
Trees_din <= "00000000011001000010110010011101";
wait for Clk_period;
Addr <= "0101011100111";
Trees_din <= "00000000000011110010110010011101";
wait for Clk_period;
Addr <= "0101011101000";
Trees_din <= "00000110000000000010011101000000";
wait for Clk_period;
Addr <= "0101011101001";
Trees_din <= "00000110000000000010000000100000";
wait for Clk_period;
Addr <= "0101011101010";
Trees_din <= "00000011000000000000101000010000";
wait for Clk_period;
Addr <= "0101011101011";
Trees_din <= "00000111000000000100001100001000";
wait for Clk_period;
Addr <= "0101011101100";
Trees_din <= "00000100000000000100000100000100";
wait for Clk_period;
Addr <= "0101011101101";
Trees_din <= "00000000001010000010110010011101";
wait for Clk_period;
Addr <= "0101011101110";
Trees_din <= "00000000001011010010110010011101";
wait for Clk_period;
Addr <= "0101011101111";
Trees_din <= "00000011000000000100010000000100";
wait for Clk_period;
Addr <= "0101011110000";
Trees_din <= "00000000001101010010110010011101";
wait for Clk_period;
Addr <= "0101011110001";
Trees_din <= "00000000001111100010110010011101";
wait for Clk_period;
Addr <= "0101011110010";
Trees_din <= "00000011000000000011100100001000";
wait for Clk_period;
Addr <= "0101011110011";
Trees_din <= "00000000000000000011101000000100";
wait for Clk_period;
Addr <= "0101011110100";
Trees_din <= "00000000010001100010110010011101";
wait for Clk_period;
Addr <= "0101011110101";
Trees_din <= "00000000000001000010110010011101";
wait for Clk_period;
Addr <= "0101011110110";
Trees_din <= "00000101000000000110000000000100";
wait for Clk_period;
Addr <= "0101011110111";
Trees_din <= "00000000010110100010110010011101";
wait for Clk_period;
Addr <= "0101011111000";
Trees_din <= "00000000010110110010110010011101";
wait for Clk_period;
Addr <= "0101011111001";
Trees_din <= "00000011000000000010100100010000";
wait for Clk_period;
Addr <= "0101011111010";
Trees_din <= "00000101000000000001111000001000";
wait for Clk_period;
Addr <= "0101011111011";
Trees_din <= "00000010000000000000110000000100";
wait for Clk_period;
Addr <= "0101011111100";
Trees_din <= "00000000011001000010110010011101";
wait for Clk_period;
Addr <= "0101011111101";
Trees_din <= "00000000010100010010110010011101";
wait for Clk_period;
Addr <= "0101011111110";
Trees_din <= "00000100000000000100000000000100";
wait for Clk_period;
Addr <= "0101011111111";
Trees_din <= "00000000010000010010110010011101";
wait for Clk_period;
Addr <= "0101100000000";
Trees_din <= "00000000011000100010110010011101";
wait for Clk_period;
Addr <= "0101100000001";
Trees_din <= "00000001000000000010111000001000";
wait for Clk_period;
Addr <= "0101100000010";
Trees_din <= "00000011000000000101101000000100";
wait for Clk_period;
Addr <= "0101100000011";
Trees_din <= "00000000000101000010110010011101";
wait for Clk_period;
Addr <= "0101100000100";
Trees_din <= "00000000010010110010110010011101";
wait for Clk_period;
Addr <= "0101100000101";
Trees_din <= "00000011000000000010100100000100";
wait for Clk_period;
Addr <= "0101100000110";
Trees_din <= "00000000000100110010110010011101";
wait for Clk_period;
Addr <= "0101100000111";
Trees_din <= "00000000000001110010110010011101";
wait for Clk_period;
Addr <= "0101100001000";
Trees_din <= "00000000000000000011001100100000";
wait for Clk_period;
Addr <= "0101100001001";
Trees_din <= "00000011000000000001101000010000";
wait for Clk_period;
Addr <= "0101100001010";
Trees_din <= "00000111000000000001001100001000";
wait for Clk_period;
Addr <= "0101100001011";
Trees_din <= "00000101000000000001000000000100";
wait for Clk_period;
Addr <= "0101100001100";
Trees_din <= "00000000000110000010110010011101";
wait for Clk_period;
Addr <= "0101100001101";
Trees_din <= "00000000010100110010110010011101";
wait for Clk_period;
Addr <= "0101100001110";
Trees_din <= "00000001000000000101111100000100";
wait for Clk_period;
Addr <= "0101100001111";
Trees_din <= "00000000000011110010110010011101";
wait for Clk_period;
Addr <= "0101100010000";
Trees_din <= "00000000000110010010110010011101";
wait for Clk_period;
Addr <= "0101100010001";
Trees_din <= "00000011000000000011011000001000";
wait for Clk_period;
Addr <= "0101100010010";
Trees_din <= "00000000000000000011101000000100";
wait for Clk_period;
Addr <= "0101100010011";
Trees_din <= "00000000000011010010110010011101";
wait for Clk_period;
Addr <= "0101100010100";
Trees_din <= "00000000010001000010110010011101";
wait for Clk_period;
Addr <= "0101100010101";
Trees_din <= "00000001000000000110010000000100";
wait for Clk_period;
Addr <= "0101100010110";
Trees_din <= "00000000000010000010110010011101";
wait for Clk_period;
Addr <= "0101100010111";
Trees_din <= "00000000010010000010110010011101";
wait for Clk_period;
Addr <= "0101100011000";
Trees_din <= "00000001000000000001011000010000";
wait for Clk_period;
Addr <= "0101100011001";
Trees_din <= "00000010000000000000000000001000";
wait for Clk_period;
Addr <= "0101100011010";
Trees_din <= "00000101000000000000000100000100";
wait for Clk_period;
Addr <= "0101100011011";
Trees_din <= "00000000000011100010110010011101";
wait for Clk_period;
Addr <= "0101100011100";
Trees_din <= "00000000001100100010110010011101";
wait for Clk_period;
Addr <= "0101100011101";
Trees_din <= "00000100000000000000110100000100";
wait for Clk_period;
Addr <= "0101100011110";
Trees_din <= "00000000010101110010110010011101";
wait for Clk_period;
Addr <= "0101100011111";
Trees_din <= "00000000000101000010110010011101";
wait for Clk_period;
Addr <= "0101100100000";
Trees_din <= "00000100000000000101000000001000";
wait for Clk_period;
Addr <= "0101100100001";
Trees_din <= "00000000000000000001111000000100";
wait for Clk_period;
Addr <= "0101100100010";
Trees_din <= "00000000011000110010110010011101";
wait for Clk_period;
Addr <= "0101100100011";
Trees_din <= "00000000000000100010110010011101";
wait for Clk_period;
Addr <= "0101100100100";
Trees_din <= "00000010000000000011111000000100";
wait for Clk_period;
Addr <= "0101100100101";
Trees_din <= "00000000010101010010110010011101";
wait for Clk_period;
Addr <= "0101100100110";
Trees_din <= "00000000001100000010110010011101";
wait for Clk_period;



----------tree 22-------------------

Addr <= "0101100100111";
Trees_din <= "00000110000000000001000110000000";
wait for Clk_period;
Addr <= "0101100101000";
Trees_din <= "00000111000000000010001101000000";
wait for Clk_period;
Addr <= "0101100101001";
Trees_din <= "00000111000000000001000100100000";
wait for Clk_period;
Addr <= "0101100101010";
Trees_din <= "00000001000000000010001000010000";
wait for Clk_period;
Addr <= "0101100101011";
Trees_din <= "00000101000000000000010100001000";
wait for Clk_period;
Addr <= "0101100101100";
Trees_din <= "00000100000000000001010100000100";
wait for Clk_period;
Addr <= "0101100101101";
Trees_din <= "00000000010110100010111010011001";
wait for Clk_period;
Addr <= "0101100101110";
Trees_din <= "00000000000101000010111010011001";
wait for Clk_period;
Addr <= "0101100101111";
Trees_din <= "00000000000000000000011100000100";
wait for Clk_period;
Addr <= "0101100110000";
Trees_din <= "00000000000111100010111010011001";
wait for Clk_period;
Addr <= "0101100110001";
Trees_din <= "00000000000010010010111010011001";
wait for Clk_period;
Addr <= "0101100110010";
Trees_din <= "00000000000000000000100100001000";
wait for Clk_period;
Addr <= "0101100110011";
Trees_din <= "00000110000000000101000000000100";
wait for Clk_period;
Addr <= "0101100110100";
Trees_din <= "00000000010100000010111010011001";
wait for Clk_period;
Addr <= "0101100110101";
Trees_din <= "00000000000101110010111010011001";
wait for Clk_period;
Addr <= "0101100110110";
Trees_din <= "00000010000000000011001100000100";
wait for Clk_period;
Addr <= "0101100110111";
Trees_din <= "00000000001000010010111010011001";
wait for Clk_period;
Addr <= "0101100111000";
Trees_din <= "00000000010101110010111010011001";
wait for Clk_period;
Addr <= "0101100111001";
Trees_din <= "00000011000000000011000100010000";
wait for Clk_period;
Addr <= "0101100111010";
Trees_din <= "00000011000000000101011000001000";
wait for Clk_period;
Addr <= "0101100111011";
Trees_din <= "00000100000000000001101100000100";
wait for Clk_period;
Addr <= "0101100111100";
Trees_din <= "00000000010110110010111010011001";
wait for Clk_period;
Addr <= "0101100111101";
Trees_din <= "00000000010011010010111010011001";
wait for Clk_period;
Addr <= "0101100111110";
Trees_din <= "00000011000000000010000000000100";
wait for Clk_period;
Addr <= "0101100111111";
Trees_din <= "00000000000000110010111010011001";
wait for Clk_period;
Addr <= "0101101000000";
Trees_din <= "00000000010110000010111010011001";
wait for Clk_period;
Addr <= "0101101000001";
Trees_din <= "00000000000000000010010000001000";
wait for Clk_period;
Addr <= "0101101000010";
Trees_din <= "00000001000000000001011100000100";
wait for Clk_period;
Addr <= "0101101000011";
Trees_din <= "00000000000101100010111010011001";
wait for Clk_period;
Addr <= "0101101000100";
Trees_din <= "00000000001101010010111010011001";
wait for Clk_period;
Addr <= "0101101000101";
Trees_din <= "00000110000000000010010000000100";
wait for Clk_period;
Addr <= "0101101000110";
Trees_din <= "00000000001010010010111010011001";
wait for Clk_period;
Addr <= "0101101000111";
Trees_din <= "00000000001110010010111010011001";
wait for Clk_period;
Addr <= "0101101001000";
Trees_din <= "00000100000000000010111000100000";
wait for Clk_period;
Addr <= "0101101001001";
Trees_din <= "00000101000000000101110000010000";
wait for Clk_period;
Addr <= "0101101001010";
Trees_din <= "00000100000000000110001000001000";
wait for Clk_period;
Addr <= "0101101001011";
Trees_din <= "00000000000000000011011100000100";
wait for Clk_period;
Addr <= "0101101001100";
Trees_din <= "00000000010010100010111010011001";
wait for Clk_period;
Addr <= "0101101001101";
Trees_din <= "00000000000110000010111010011001";
wait for Clk_period;
Addr <= "0101101001110";
Trees_din <= "00000101000000000110000000000100";
wait for Clk_period;
Addr <= "0101101001111";
Trees_din <= "00000000000101000010111010011001";
wait for Clk_period;
Addr <= "0101101010000";
Trees_din <= "00000000000101010010111010011001";
wait for Clk_period;
Addr <= "0101101010001";
Trees_din <= "00000001000000000100110000001000";
wait for Clk_period;
Addr <= "0101101010010";
Trees_din <= "00000011000000000100000100000100";
wait for Clk_period;
Addr <= "0101101010011";
Trees_din <= "00000000001100110010111010011001";
wait for Clk_period;
Addr <= "0101101010100";
Trees_din <= "00000000000010010010111010011001";
wait for Clk_period;
Addr <= "0101101010101";
Trees_din <= "00000011000000000101010000000100";
wait for Clk_period;
Addr <= "0101101010110";
Trees_din <= "00000000001101010010111010011001";
wait for Clk_period;
Addr <= "0101101010111";
Trees_din <= "00000000000110100010111010011001";
wait for Clk_period;
Addr <= "0101101011000";
Trees_din <= "00000010000000000100011000010000";
wait for Clk_period;
Addr <= "0101101011001";
Trees_din <= "00000010000000000000001000001000";
wait for Clk_period;
Addr <= "0101101011010";
Trees_din <= "00000101000000000101001100000100";
wait for Clk_period;
Addr <= "0101101011011";
Trees_din <= "00000000001000100010111010011001";
wait for Clk_period;
Addr <= "0101101011100";
Trees_din <= "00000000001100110010111010011001";
wait for Clk_period;
Addr <= "0101101011101";
Trees_din <= "00000100000000000011111100000100";
wait for Clk_period;
Addr <= "0101101011110";
Trees_din <= "00000000010110000010111010011001";
wait for Clk_period;
Addr <= "0101101011111";
Trees_din <= "00000000010111000010111010011001";
wait for Clk_period;
Addr <= "0101101100000";
Trees_din <= "00000000000000000010111100001000";
wait for Clk_period;
Addr <= "0101101100001";
Trees_din <= "00000110000000000011000000000100";
wait for Clk_period;
Addr <= "0101101100010";
Trees_din <= "00000000000100000010111010011001";
wait for Clk_period;
Addr <= "0101101100011";
Trees_din <= "00000000001110000010111010011001";
wait for Clk_period;
Addr <= "0101101100100";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "0101101100101";
Trees_din <= "00000000010001010010111010011001";
wait for Clk_period;
Addr <= "0101101100110";
Trees_din <= "00000000000110000010111010011001";
wait for Clk_period;
Addr <= "0101101100111";
Trees_din <= "00000011000000000001111001000000";
wait for Clk_period;
Addr <= "0101101101000";
Trees_din <= "00000110000000000101101000100000";
wait for Clk_period;
Addr <= "0101101101001";
Trees_din <= "00000110000000000101000100010000";
wait for Clk_period;
Addr <= "0101101101010";
Trees_din <= "00000100000000000101001100001000";
wait for Clk_period;
Addr <= "0101101101011";
Trees_din <= "00000100000000000101110100000100";
wait for Clk_period;
Addr <= "0101101101100";
Trees_din <= "00000000000001100010111010011001";
wait for Clk_period;
Addr <= "0101101101101";
Trees_din <= "00000000010001110010111010011001";
wait for Clk_period;
Addr <= "0101101101110";
Trees_din <= "00000011000000000001000000000100";
wait for Clk_period;
Addr <= "0101101101111";
Trees_din <= "00000000000101100010111010011001";
wait for Clk_period;
Addr <= "0101101110000";
Trees_din <= "00000000000011000010111010011001";
wait for Clk_period;
Addr <= "0101101110001";
Trees_din <= "00000111000000000000110100001000";
wait for Clk_period;
Addr <= "0101101110010";
Trees_din <= "00000111000000000100010000000100";
wait for Clk_period;
Addr <= "0101101110011";
Trees_din <= "00000000001110010010111010011001";
wait for Clk_period;
Addr <= "0101101110100";
Trees_din <= "00000000000011010010111010011001";
wait for Clk_period;
Addr <= "0101101110101";
Trees_din <= "00000011000000000011101000000100";
wait for Clk_period;
Addr <= "0101101110110";
Trees_din <= "00000000001010010010111010011001";
wait for Clk_period;
Addr <= "0101101110111";
Trees_din <= "00000000001100010010111010011001";
wait for Clk_period;
Addr <= "0101101111000";
Trees_din <= "00000011000000000011000100010000";
wait for Clk_period;
Addr <= "0101101111001";
Trees_din <= "00000100000000000100100000001000";
wait for Clk_period;
Addr <= "0101101111010";
Trees_din <= "00000111000000000001100000000100";
wait for Clk_period;
Addr <= "0101101111011";
Trees_din <= "00000000010110000010111010011001";
wait for Clk_period;
Addr <= "0101101111100";
Trees_din <= "00000000010110110010111010011001";
wait for Clk_period;
Addr <= "0101101111101";
Trees_din <= "00000010000000000001100100000100";
wait for Clk_period;
Addr <= "0101101111110";
Trees_din <= "00000000001101010010111010011001";
wait for Clk_period;
Addr <= "0101101111111";
Trees_din <= "00000000011000110010111010011001";
wait for Clk_period;
Addr <= "0101110000000";
Trees_din <= "00000101000000000100011000001000";
wait for Clk_period;
Addr <= "0101110000001";
Trees_din <= "00000001000000000101111000000100";
wait for Clk_period;
Addr <= "0101110000010";
Trees_din <= "00000000001010010010111010011001";
wait for Clk_period;
Addr <= "0101110000011";
Trees_din <= "00000000010110010010111010011001";
wait for Clk_period;
Addr <= "0101110000100";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "0101110000101";
Trees_din <= "00000000011000110010111010011001";
wait for Clk_period;
Addr <= "0101110000110";
Trees_din <= "00000000010011000010111010011001";
wait for Clk_period;
Addr <= "0101110000111";
Trees_din <= "00000110000000000001011000100000";
wait for Clk_period;
Addr <= "0101110001000";
Trees_din <= "00000111000000000101110100010000";
wait for Clk_period;
Addr <= "0101110001001";
Trees_din <= "00000000000000000011011100001000";
wait for Clk_period;
Addr <= "0101110001010";
Trees_din <= "00000001000000000100100100000100";
wait for Clk_period;
Addr <= "0101110001011";
Trees_din <= "00000000010011100010111010011001";
wait for Clk_period;
Addr <= "0101110001100";
Trees_din <= "00000000001101010010111010011001";
wait for Clk_period;
Addr <= "0101110001101";
Trees_din <= "00000101000000000101001000000100";
wait for Clk_period;
Addr <= "0101110001110";
Trees_din <= "00000000000110010010111010011001";
wait for Clk_period;
Addr <= "0101110001111";
Trees_din <= "00000000000111000010111010011001";
wait for Clk_period;
Addr <= "0101110010000";
Trees_din <= "00000111000000000000011100001000";
wait for Clk_period;
Addr <= "0101110010001";
Trees_din <= "00000101000000000101011100000100";
wait for Clk_period;
Addr <= "0101110010010";
Trees_din <= "00000000010111010010111010011001";
wait for Clk_period;
Addr <= "0101110010011";
Trees_din <= "00000000000111010010111010011001";
wait for Clk_period;
Addr <= "0101110010100";
Trees_din <= "00000101000000000100101100000100";
wait for Clk_period;
Addr <= "0101110010101";
Trees_din <= "00000000010010010010111010011001";
wait for Clk_period;
Addr <= "0101110010110";
Trees_din <= "00000000000100010010111010011001";
wait for Clk_period;
Addr <= "0101110010111";
Trees_din <= "00000001000000000100001100010000";
wait for Clk_period;
Addr <= "0101110011000";
Trees_din <= "00000000000000000011011000001000";
wait for Clk_period;
Addr <= "0101110011001";
Trees_din <= "00000001000000000011110100000100";
wait for Clk_period;
Addr <= "0101110011010";
Trees_din <= "00000000001110000010111010011001";
wait for Clk_period;
Addr <= "0101110011011";
Trees_din <= "00000000010110010010111010011001";
wait for Clk_period;
Addr <= "0101110011100";
Trees_din <= "00000010000000000011111100000100";
wait for Clk_period;
Addr <= "0101110011101";
Trees_din <= "00000000010101010010111010011001";
wait for Clk_period;
Addr <= "0101110011110";
Trees_din <= "00000000010111100010111010011001";
wait for Clk_period;
Addr <= "0101110011111";
Trees_din <= "00000100000000000101011000001000";
wait for Clk_period;
Addr <= "0101110100000";
Trees_din <= "00000110000000000010101100000100";
wait for Clk_period;
Addr <= "0101110100001";
Trees_din <= "00000000010111000010111010011001";
wait for Clk_period;
Addr <= "0101110100010";
Trees_din <= "00000000011000110010111010011001";
wait for Clk_period;
Addr <= "0101110100011";
Trees_din <= "00000011000000000010100000000100";
wait for Clk_period;
Addr <= "0101110100100";
Trees_din <= "00000000000001110010111010011001";
wait for Clk_period;
Addr <= "0101110100101";
Trees_din <= "00000000000001000010111010011001";
wait for Clk_period;



----------tree 23-------------------

Addr <= "0101110100110";
Trees_din <= "00000111000000000011011110000000";
wait for Clk_period;
Addr <= "0101110100111";
Trees_din <= "00000111000000000010111101000000";
wait for Clk_period;
Addr <= "0101110101000";
Trees_din <= "00000011000000000010111000100000";
wait for Clk_period;
Addr <= "0101110101001";
Trees_din <= "00000001000000000010111100010000";
wait for Clk_period;
Addr <= "0101110101010";
Trees_din <= "00000011000000000000001100001000";
wait for Clk_period;
Addr <= "0101110101011";
Trees_din <= "00000110000000000010000100000100";
wait for Clk_period;
Addr <= "0101110101100";
Trees_din <= "00000000010010010011000010010101";
wait for Clk_period;
Addr <= "0101110101101";
Trees_din <= "00000000000001110011000010010101";
wait for Clk_period;
Addr <= "0101110101110";
Trees_din <= "00000110000000000000100000000100";
wait for Clk_period;
Addr <= "0101110101111";
Trees_din <= "00000000000111000011000010010101";
wait for Clk_period;
Addr <= "0101110110000";
Trees_din <= "00000000000110000011000010010101";
wait for Clk_period;
Addr <= "0101110110001";
Trees_din <= "00000001000000000011001100001000";
wait for Clk_period;
Addr <= "0101110110010";
Trees_din <= "00000010000000000000000000000100";
wait for Clk_period;
Addr <= "0101110110011";
Trees_din <= "00000000010110100011000010010101";
wait for Clk_period;
Addr <= "0101110110100";
Trees_din <= "00000000001110110011000010010101";
wait for Clk_period;
Addr <= "0101110110101";
Trees_din <= "00000011000000000100001100000100";
wait for Clk_period;
Addr <= "0101110110110";
Trees_din <= "00000000000100100011000010010101";
wait for Clk_period;
Addr <= "0101110110111";
Trees_din <= "00000000000001000011000010010101";
wait for Clk_period;
Addr <= "0101110111000";
Trees_din <= "00000011000000000010011000010000";
wait for Clk_period;
Addr <= "0101110111001";
Trees_din <= "00000100000000000001110100001000";
wait for Clk_period;
Addr <= "0101110111010";
Trees_din <= "00000111000000000010101000000100";
wait for Clk_period;
Addr <= "0101110111011";
Trees_din <= "00000000011000010011000010010101";
wait for Clk_period;
Addr <= "0101110111100";
Trees_din <= "00000000001001100011000010010101";
wait for Clk_period;
Addr <= "0101110111101";
Trees_din <= "00000100000000000110001100000100";
wait for Clk_period;
Addr <= "0101110111110";
Trees_din <= "00000000010111110011000010010101";
wait for Clk_period;
Addr <= "0101110111111";
Trees_din <= "00000000000000010011000010010101";
wait for Clk_period;
Addr <= "0101111000000";
Trees_din <= "00000101000000000000011000001000";
wait for Clk_period;
Addr <= "0101111000001";
Trees_din <= "00000100000000000000011000000100";
wait for Clk_period;
Addr <= "0101111000010";
Trees_din <= "00000000011000000011000010010101";
wait for Clk_period;
Addr <= "0101111000011";
Trees_din <= "00000000001101000011000010010101";
wait for Clk_period;
Addr <= "0101111000100";
Trees_din <= "00000000000000000010101000000100";
wait for Clk_period;
Addr <= "0101111000101";
Trees_din <= "00000000000000100011000010010101";
wait for Clk_period;
Addr <= "0101111000110";
Trees_din <= "00000000001110000011000010010101";
wait for Clk_period;
Addr <= "0101111000111";
Trees_din <= "00000101000000000100010000100000";
wait for Clk_period;
Addr <= "0101111001000";
Trees_din <= "00000101000000000000011000010000";
wait for Clk_period;
Addr <= "0101111001001";
Trees_din <= "00000100000000000001011100001000";
wait for Clk_period;
Addr <= "0101111001010";
Trees_din <= "00000101000000000001011100000100";
wait for Clk_period;
Addr <= "0101111001011";
Trees_din <= "00000000000001110011000010010101";
wait for Clk_period;
Addr <= "0101111001100";
Trees_din <= "00000000011000100011000010010101";
wait for Clk_period;
Addr <= "0101111001101";
Trees_din <= "00000111000000000001010000000100";
wait for Clk_period;
Addr <= "0101111001110";
Trees_din <= "00000000000011100011000010010101";
wait for Clk_period;
Addr <= "0101111001111";
Trees_din <= "00000000000111000011000010010101";
wait for Clk_period;
Addr <= "0101111010000";
Trees_din <= "00000111000000000101000000001000";
wait for Clk_period;
Addr <= "0101111010001";
Trees_din <= "00000111000000000101001100000100";
wait for Clk_period;
Addr <= "0101111010010";
Trees_din <= "00000000000001010011000010010101";
wait for Clk_period;
Addr <= "0101111010011";
Trees_din <= "00000000000001110011000010010101";
wait for Clk_period;
Addr <= "0101111010100";
Trees_din <= "00000101000000000100011100000100";
wait for Clk_period;
Addr <= "0101111010101";
Trees_din <= "00000000000010100011000010010101";
wait for Clk_period;
Addr <= "0101111010110";
Trees_din <= "00000000001111010011000010010101";
wait for Clk_period;
Addr <= "0101111010111";
Trees_din <= "00000010000000000010111000010000";
wait for Clk_period;
Addr <= "0101111011000";
Trees_din <= "00000000000000000101000100001000";
wait for Clk_period;
Addr <= "0101111011001";
Trees_din <= "00000011000000000001100000000100";
wait for Clk_period;
Addr <= "0101111011010";
Trees_din <= "00000000000000000011000010010101";
wait for Clk_period;
Addr <= "0101111011011";
Trees_din <= "00000000001100010011000010010101";
wait for Clk_period;
Addr <= "0101111011100";
Trees_din <= "00000010000000000010111000000100";
wait for Clk_period;
Addr <= "0101111011101";
Trees_din <= "00000000001000110011000010010101";
wait for Clk_period;
Addr <= "0101111011110";
Trees_din <= "00000000001000010011000010010101";
wait for Clk_period;
Addr <= "0101111011111";
Trees_din <= "00000100000000000000000100001000";
wait for Clk_period;
Addr <= "0101111100000";
Trees_din <= "00000111000000000000111000000100";
wait for Clk_period;
Addr <= "0101111100001";
Trees_din <= "00000000000010010011000010010101";
wait for Clk_period;
Addr <= "0101111100010";
Trees_din <= "00000000000011100011000010010101";
wait for Clk_period;
Addr <= "0101111100011";
Trees_din <= "00000011000000000000100000000100";
wait for Clk_period;
Addr <= "0101111100100";
Trees_din <= "00000000001100100011000010010101";
wait for Clk_period;
Addr <= "0101111100101";
Trees_din <= "00000000000000010011000010010101";
wait for Clk_period;
Addr <= "0101111100110";
Trees_din <= "00000100000000000010001101000000";
wait for Clk_period;
Addr <= "0101111100111";
Trees_din <= "00000110000000000100010100100000";
wait for Clk_period;
Addr <= "0101111101000";
Trees_din <= "00000010000000000001100000010000";
wait for Clk_period;
Addr <= "0101111101001";
Trees_din <= "00000111000000000011101000001000";
wait for Clk_period;
Addr <= "0101111101010";
Trees_din <= "00000101000000000011010100000100";
wait for Clk_period;
Addr <= "0101111101011";
Trees_din <= "00000000001111100011000010010101";
wait for Clk_period;
Addr <= "0101111101100";
Trees_din <= "00000000000100100011000010010101";
wait for Clk_period;
Addr <= "0101111101101";
Trees_din <= "00000111000000000010001100000100";
wait for Clk_period;
Addr <= "0101111101110";
Trees_din <= "00000000000010000011000010010101";
wait for Clk_period;
Addr <= "0101111101111";
Trees_din <= "00000000000100110011000010010101";
wait for Clk_period;
Addr <= "0101111110000";
Trees_din <= "00000010000000000101001100001000";
wait for Clk_period;
Addr <= "0101111110001";
Trees_din <= "00000000000000000110001000000100";
wait for Clk_period;
Addr <= "0101111110010";
Trees_din <= "00000000010110110011000010010101";
wait for Clk_period;
Addr <= "0101111110011";
Trees_din <= "00000000010001110011000010010101";
wait for Clk_period;
Addr <= "0101111110100";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "0101111110101";
Trees_din <= "00000000010100010011000010010101";
wait for Clk_period;
Addr <= "0101111110110";
Trees_din <= "00000000010101000011000010010101";
wait for Clk_period;
Addr <= "0101111110111";
Trees_din <= "00000011000000000100110100010000";
wait for Clk_period;
Addr <= "0101111111000";
Trees_din <= "00000101000000000001100100001000";
wait for Clk_period;
Addr <= "0101111111001";
Trees_din <= "00000000000000000010000000000100";
wait for Clk_period;
Addr <= "0101111111010";
Trees_din <= "00000000010101100011000010010101";
wait for Clk_period;
Addr <= "0101111111011";
Trees_din <= "00000000001011110011000010010101";
wait for Clk_period;
Addr <= "0101111111100";
Trees_din <= "00000010000000000101010000000100";
wait for Clk_period;
Addr <= "0101111111101";
Trees_din <= "00000000010101100011000010010101";
wait for Clk_period;
Addr <= "0101111111110";
Trees_din <= "00000000010001100011000010010101";
wait for Clk_period;
Addr <= "0101111111111";
Trees_din <= "00000000000000000010000000001000";
wait for Clk_period;
Addr <= "0110000000000";
Trees_din <= "00000001000000000001000100000100";
wait for Clk_period;
Addr <= "0110000000001";
Trees_din <= "00000000001011110011000010010101";
wait for Clk_period;
Addr <= "0110000000010";
Trees_din <= "00000000011000110011000010010101";
wait for Clk_period;
Addr <= "0110000000011";
Trees_din <= "00000001000000000101111000000100";
wait for Clk_period;
Addr <= "0110000000100";
Trees_din <= "00000000000010000011000010010101";
wait for Clk_period;
Addr <= "0110000000101";
Trees_din <= "00000000011000000011000010010101";
wait for Clk_period;
Addr <= "0110000000110";
Trees_din <= "00000110000000000011010100100000";
wait for Clk_period;
Addr <= "0110000000111";
Trees_din <= "00000011000000000000000100010000";
wait for Clk_period;
Addr <= "0110000001000";
Trees_din <= "00000001000000000100100100001000";
wait for Clk_period;
Addr <= "0110000001001";
Trees_din <= "00000111000000000001100000000100";
wait for Clk_period;
Addr <= "0110000001010";
Trees_din <= "00000000001001000011000010010101";
wait for Clk_period;
Addr <= "0110000001011";
Trees_din <= "00000000000011110011000010010101";
wait for Clk_period;
Addr <= "0110000001100";
Trees_din <= "00000100000000000101110100000100";
wait for Clk_period;
Addr <= "0110000001101";
Trees_din <= "00000000000111100011000010010101";
wait for Clk_period;
Addr <= "0110000001110";
Trees_din <= "00000000001111110011000010010101";
wait for Clk_period;
Addr <= "0110000001111";
Trees_din <= "00000100000000000100010000001000";
wait for Clk_period;
Addr <= "0110000010000";
Trees_din <= "00000101000000000011100000000100";
wait for Clk_period;
Addr <= "0110000010001";
Trees_din <= "00000000010000010011000010010101";
wait for Clk_period;
Addr <= "0110000010010";
Trees_din <= "00000000000100100011000010010101";
wait for Clk_period;
Addr <= "0110000010011";
Trees_din <= "00000000000000000101101100000100";
wait for Clk_period;
Addr <= "0110000010100";
Trees_din <= "00000000001101010011000010010101";
wait for Clk_period;
Addr <= "0110000010101";
Trees_din <= "00000000000111110011000010010101";
wait for Clk_period;
Addr <= "0110000010110";
Trees_din <= "00000100000000000100110000010000";
wait for Clk_period;
Addr <= "0110000010111";
Trees_din <= "00000110000000000000101100001000";
wait for Clk_period;
Addr <= "0110000011000";
Trees_din <= "00000101000000000011110000000100";
wait for Clk_period;
Addr <= "0110000011001";
Trees_din <= "00000000010111110011000010010101";
wait for Clk_period;
Addr <= "0110000011010";
Trees_din <= "00000000001110000011000010010101";
wait for Clk_period;
Addr <= "0110000011011";
Trees_din <= "00000011000000000010001000000100";
wait for Clk_period;
Addr <= "0110000011100";
Trees_din <= "00000000001011110011000010010101";
wait for Clk_period;
Addr <= "0110000011101";
Trees_din <= "00000000000100110011000010010101";
wait for Clk_period;
Addr <= "0110000011110";
Trees_din <= "00000010000000000101011000001000";
wait for Clk_period;
Addr <= "0110000011111";
Trees_din <= "00000011000000000110001100000100";
wait for Clk_period;
Addr <= "0110000100000";
Trees_din <= "00000000001111010011000010010101";
wait for Clk_period;
Addr <= "0110000100001";
Trees_din <= "00000000011000000011000010010101";
wait for Clk_period;
Addr <= "0110000100010";
Trees_din <= "00000000000000000010011100000100";
wait for Clk_period;
Addr <= "0110000100011";
Trees_din <= "00000000001100110011000010010101";
wait for Clk_period;
Addr <= "0110000100100";
Trees_din <= "00000000001001010011000010010101";
wait for Clk_period;



----------tree 24-------------------

Addr <= "0110000100101";
Trees_din <= "00000001000000000001010010000000";
wait for Clk_period;
Addr <= "0110000100110";
Trees_din <= "00000001000000000010010101000000";
wait for Clk_period;
Addr <= "0110000100111";
Trees_din <= "00000010000000000100001100100000";
wait for Clk_period;
Addr <= "0110000101000";
Trees_din <= "00000101000000000000001000010000";
wait for Clk_period;
Addr <= "0110000101001";
Trees_din <= "00000101000000000011100000001000";
wait for Clk_period;
Addr <= "0110000101010";
Trees_din <= "00000010000000000101010100000100";
wait for Clk_period;
Addr <= "0110000101011";
Trees_din <= "00000000000110000011001010010001";
wait for Clk_period;
Addr <= "0110000101100";
Trees_din <= "00000000001011000011001010010001";
wait for Clk_period;
Addr <= "0110000101101";
Trees_din <= "00000010000000000100100000000100";
wait for Clk_period;
Addr <= "0110000101110";
Trees_din <= "00000000011000010011001010010001";
wait for Clk_period;
Addr <= "0110000101111";
Trees_din <= "00000000000101000011001010010001";
wait for Clk_period;
Addr <= "0110000110000";
Trees_din <= "00000000000000000011100000001000";
wait for Clk_period;
Addr <= "0110000110001";
Trees_din <= "00000110000000000000111000000100";
wait for Clk_period;
Addr <= "0110000110010";
Trees_din <= "00000000010110010011001010010001";
wait for Clk_period;
Addr <= "0110000110011";
Trees_din <= "00000000001101100011001010010001";
wait for Clk_period;
Addr <= "0110000110100";
Trees_din <= "00000110000000000000000000000100";
wait for Clk_period;
Addr <= "0110000110101";
Trees_din <= "00000000000110110011001010010001";
wait for Clk_period;
Addr <= "0110000110110";
Trees_din <= "00000000000101100011001010010001";
wait for Clk_period;
Addr <= "0110000110111";
Trees_din <= "00000101000000000000101000010000";
wait for Clk_period;
Addr <= "0110000111000";
Trees_din <= "00000111000000000001011100001000";
wait for Clk_period;
Addr <= "0110000111001";
Trees_din <= "00000000000000000001111000000100";
wait for Clk_period;
Addr <= "0110000111010";
Trees_din <= "00000000010100010011001010010001";
wait for Clk_period;
Addr <= "0110000111011";
Trees_din <= "00000000000011100011001010010001";
wait for Clk_period;
Addr <= "0110000111100";
Trees_din <= "00000101000000000001010000000100";
wait for Clk_period;
Addr <= "0110000111101";
Trees_din <= "00000000000011010011001010010001";
wait for Clk_period;
Addr <= "0110000111110";
Trees_din <= "00000000001000100011001010010001";
wait for Clk_period;
Addr <= "0110000111111";
Trees_din <= "00000100000000000010001000001000";
wait for Clk_period;
Addr <= "0110001000000";
Trees_din <= "00000010000000000101010000000100";
wait for Clk_period;
Addr <= "0110001000001";
Trees_din <= "00000000000110000011001010010001";
wait for Clk_period;
Addr <= "0110001000010";
Trees_din <= "00000000000111110011001010010001";
wait for Clk_period;
Addr <= "0110001000011";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "0110001000100";
Trees_din <= "00000000001110000011001010010001";
wait for Clk_period;
Addr <= "0110001000101";
Trees_din <= "00000000001110100011001010010001";
wait for Clk_period;
Addr <= "0110001000110";
Trees_din <= "00000101000000000100011100100000";
wait for Clk_period;
Addr <= "0110001000111";
Trees_din <= "00000101000000000001010000010000";
wait for Clk_period;
Addr <= "0110001001000";
Trees_din <= "00000111000000000000010000001000";
wait for Clk_period;
Addr <= "0110001001001";
Trees_din <= "00000001000000000010011000000100";
wait for Clk_period;
Addr <= "0110001001010";
Trees_din <= "00000000010011010011001010010001";
wait for Clk_period;
Addr <= "0110001001011";
Trees_din <= "00000000010000000011001010010001";
wait for Clk_period;
Addr <= "0110001001100";
Trees_din <= "00000001000000000101110000000100";
wait for Clk_period;
Addr <= "0110001001101";
Trees_din <= "00000000001001010011001010010001";
wait for Clk_period;
Addr <= "0110001001110";
Trees_din <= "00000000011001000011001010010001";
wait for Clk_period;
Addr <= "0110001001111";
Trees_din <= "00000001000000000001011100001000";
wait for Clk_period;
Addr <= "0110001010000";
Trees_din <= "00000010000000000011010000000100";
wait for Clk_period;
Addr <= "0110001010001";
Trees_din <= "00000000000000110011001010010001";
wait for Clk_period;
Addr <= "0110001010010";
Trees_din <= "00000000000010000011001010010001";
wait for Clk_period;
Addr <= "0110001010011";
Trees_din <= "00000000000000000100000100000100";
wait for Clk_period;
Addr <= "0110001010100";
Trees_din <= "00000000000000110011001010010001";
wait for Clk_period;
Addr <= "0110001010101";
Trees_din <= "00000000000001000011001010010001";
wait for Clk_period;
Addr <= "0110001010110";
Trees_din <= "00000110000000000100110000010000";
wait for Clk_period;
Addr <= "0110001010111";
Trees_din <= "00000000000000000001011000001000";
wait for Clk_period;
Addr <= "0110001011000";
Trees_din <= "00000100000000000100100100000100";
wait for Clk_period;
Addr <= "0110001011001";
Trees_din <= "00000000001001100011001010010001";
wait for Clk_period;
Addr <= "0110001011010";
Trees_din <= "00000000000011010011001010010001";
wait for Clk_period;
Addr <= "0110001011011";
Trees_din <= "00000101000000000101001100000100";
wait for Clk_period;
Addr <= "0110001011100";
Trees_din <= "00000000010000010011001010010001";
wait for Clk_period;
Addr <= "0110001011101";
Trees_din <= "00000000000001000011001010010001";
wait for Clk_period;
Addr <= "0110001011110";
Trees_din <= "00000010000000000100000000001000";
wait for Clk_period;
Addr <= "0110001011111";
Trees_din <= "00000110000000000001011000000100";
wait for Clk_period;
Addr <= "0110001100000";
Trees_din <= "00000000010010000011001010010001";
wait for Clk_period;
Addr <= "0110001100001";
Trees_din <= "00000000001111100011001010010001";
wait for Clk_period;
Addr <= "0110001100010";
Trees_din <= "00000110000000000000101000000100";
wait for Clk_period;
Addr <= "0110001100011";
Trees_din <= "00000000000010010011001010010001";
wait for Clk_period;
Addr <= "0110001100100";
Trees_din <= "00000000010100000011001010010001";
wait for Clk_period;
Addr <= "0110001100101";
Trees_din <= "00000111000000000100001001000000";
wait for Clk_period;
Addr <= "0110001100110";
Trees_din <= "00000001000000000010011100100000";
wait for Clk_period;
Addr <= "0110001100111";
Trees_din <= "00000001000000000100100000010000";
wait for Clk_period;
Addr <= "0110001101000";
Trees_din <= "00000010000000000011100100001000";
wait for Clk_period;
Addr <= "0110001101001";
Trees_din <= "00000010000000000010010000000100";
wait for Clk_period;
Addr <= "0110001101010";
Trees_din <= "00000000010000000011001010010001";
wait for Clk_period;
Addr <= "0110001101011";
Trees_din <= "00000000001101010011001010010001";
wait for Clk_period;
Addr <= "0110001101100";
Trees_din <= "00000111000000000010101100000100";
wait for Clk_period;
Addr <= "0110001101101";
Trees_din <= "00000000000111010011001010010001";
wait for Clk_period;
Addr <= "0110001101110";
Trees_din <= "00000000010100100011001010010001";
wait for Clk_period;
Addr <= "0110001101111";
Trees_din <= "00000101000000000011011100001000";
wait for Clk_period;
Addr <= "0110001110000";
Trees_din <= "00000100000000000100111000000100";
wait for Clk_period;
Addr <= "0110001110001";
Trees_din <= "00000000010101110011001010010001";
wait for Clk_period;
Addr <= "0110001110010";
Trees_din <= "00000000000001110011001010010001";
wait for Clk_period;
Addr <= "0110001110011";
Trees_din <= "00000110000000000110001100000100";
wait for Clk_period;
Addr <= "0110001110100";
Trees_din <= "00000000000101110011001010010001";
wait for Clk_period;
Addr <= "0110001110101";
Trees_din <= "00000000000001100011001010010001";
wait for Clk_period;
Addr <= "0110001110110";
Trees_din <= "00000110000000000100000000010000";
wait for Clk_period;
Addr <= "0110001110111";
Trees_din <= "00000111000000000000110000001000";
wait for Clk_period;
Addr <= "0110001111000";
Trees_din <= "00000001000000000001100100000100";
wait for Clk_period;
Addr <= "0110001111001";
Trees_din <= "00000000000101110011001010010001";
wait for Clk_period;
Addr <= "0110001111010";
Trees_din <= "00000000011000010011001010010001";
wait for Clk_period;
Addr <= "0110001111011";
Trees_din <= "00000110000000000101000100000100";
wait for Clk_period;
Addr <= "0110001111100";
Trees_din <= "00000000010010110011001010010001";
wait for Clk_period;
Addr <= "0110001111101";
Trees_din <= "00000000001110100011001010010001";
wait for Clk_period;
Addr <= "0110001111110";
Trees_din <= "00000011000000000001000100001000";
wait for Clk_period;
Addr <= "0110001111111";
Trees_din <= "00000010000000000000110000000100";
wait for Clk_period;
Addr <= "0110010000000";
Trees_din <= "00000000001110110011001010010001";
wait for Clk_period;
Addr <= "0110010000001";
Trees_din <= "00000000010010000011001010010001";
wait for Clk_period;
Addr <= "0110010000010";
Trees_din <= "00000111000000000101111000000100";
wait for Clk_period;
Addr <= "0110010000011";
Trees_din <= "00000000001101010011001010010001";
wait for Clk_period;
Addr <= "0110010000100";
Trees_din <= "00000000001101110011001010010001";
wait for Clk_period;
Addr <= "0110010000101";
Trees_din <= "00000001000000000101001000100000";
wait for Clk_period;
Addr <= "0110010000110";
Trees_din <= "00000110000000000010101000010000";
wait for Clk_period;
Addr <= "0110010000111";
Trees_din <= "00000010000000000001100100001000";
wait for Clk_period;
Addr <= "0110010001000";
Trees_din <= "00000000000000000101011100000100";
wait for Clk_period;
Addr <= "0110010001001";
Trees_din <= "00000000000110110011001010010001";
wait for Clk_period;
Addr <= "0110010001010";
Trees_din <= "00000000000000010011001010010001";
wait for Clk_period;
Addr <= "0110010001011";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "0110010001100";
Trees_din <= "00000000010100000011001010010001";
wait for Clk_period;
Addr <= "0110010001101";
Trees_din <= "00000000001011000011001010010001";
wait for Clk_period;
Addr <= "0110010001110";
Trees_din <= "00000000000000000010011000001000";
wait for Clk_period;
Addr <= "0110010001111";
Trees_din <= "00000101000000000000101100000100";
wait for Clk_period;
Addr <= "0110010010000";
Trees_din <= "00000000001100010011001010010001";
wait for Clk_period;
Addr <= "0110010010001";
Trees_din <= "00000000010110100011001010010001";
wait for Clk_period;
Addr <= "0110010010010";
Trees_din <= "00000111000000000011010100000100";
wait for Clk_period;
Addr <= "0110010010011";
Trees_din <= "00000000010101110011001010010001";
wait for Clk_period;
Addr <= "0110010010100";
Trees_din <= "00000000001101010011001010010001";
wait for Clk_period;
Addr <= "0110010010101";
Trees_din <= "00000010000000000011111100010000";
wait for Clk_period;
Addr <= "0110010010110";
Trees_din <= "00000101000000000000010100001000";
wait for Clk_period;
Addr <= "0110010010111";
Trees_din <= "00000110000000000000010000000100";
wait for Clk_period;
Addr <= "0110010011000";
Trees_din <= "00000000000100010011001010010001";
wait for Clk_period;
Addr <= "0110010011001";
Trees_din <= "00000000000010100011001010010001";
wait for Clk_period;
Addr <= "0110010011010";
Trees_din <= "00000111000000000010111000000100";
wait for Clk_period;
Addr <= "0110010011011";
Trees_din <= "00000000010111010011001010010001";
wait for Clk_period;
Addr <= "0110010011100";
Trees_din <= "00000000000010110011001010010001";
wait for Clk_period;
Addr <= "0110010011101";
Trees_din <= "00000011000000000000001000001000";
wait for Clk_period;
Addr <= "0110010011110";
Trees_din <= "00000000000000000001011000000100";
wait for Clk_period;
Addr <= "0110010011111";
Trees_din <= "00000000001011110011001010010001";
wait for Clk_period;
Addr <= "0110010100000";
Trees_din <= "00000000001011010011001010010001";
wait for Clk_period;
Addr <= "0110010100001";
Trees_din <= "00000010000000000011011000000100";
wait for Clk_period;
Addr <= "0110010100010";
Trees_din <= "00000000000011110011001010010001";
wait for Clk_period;
Addr <= "0110010100011";
Trees_din <= "00000000000101100011001010010001";
wait for Clk_period;



----------tree 25-------------------

Addr <= "0110010100100";
Trees_din <= "00000110000000000011001010000000";
wait for Clk_period;
Addr <= "0110010100101";
Trees_din <= "00000000000000000001000101000000";
wait for Clk_period;
Addr <= "0110010100110";
Trees_din <= "00000100000000000000000100100000";
wait for Clk_period;
Addr <= "0110010100111";
Trees_din <= "00000000000000000101110100010000";
wait for Clk_period;
Addr <= "0110010101000";
Trees_din <= "00000000000000000010111000001000";
wait for Clk_period;
Addr <= "0110010101001";
Trees_din <= "00000100000000000010010000000100";
wait for Clk_period;
Addr <= "0110010101010";
Trees_din <= "00000000010111010011010010001101";
wait for Clk_period;
Addr <= "0110010101011";
Trees_din <= "00000000000001000011010010001101";
wait for Clk_period;
Addr <= "0110010101100";
Trees_din <= "00000000000000000000001000000100";
wait for Clk_period;
Addr <= "0110010101101";
Trees_din <= "00000000001000110011010010001101";
wait for Clk_period;
Addr <= "0110010101110";
Trees_din <= "00000000000111100011010010001101";
wait for Clk_period;
Addr <= "0110010101111";
Trees_din <= "00000011000000000100110100001000";
wait for Clk_period;
Addr <= "0110010110000";
Trees_din <= "00000111000000000101001100000100";
wait for Clk_period;
Addr <= "0110010110001";
Trees_din <= "00000000010110100011010010001101";
wait for Clk_period;
Addr <= "0110010110010";
Trees_din <= "00000000000101010011010010001101";
wait for Clk_period;
Addr <= "0110010110011";
Trees_din <= "00000111000000000001111100000100";
wait for Clk_period;
Addr <= "0110010110100";
Trees_din <= "00000000001101100011010010001101";
wait for Clk_period;
Addr <= "0110010110101";
Trees_din <= "00000000001010110011010010001101";
wait for Clk_period;
Addr <= "0110010110110";
Trees_din <= "00000010000000000100010000010000";
wait for Clk_period;
Addr <= "0110010110111";
Trees_din <= "00000000000000000000100000001000";
wait for Clk_period;
Addr <= "0110010111000";
Trees_din <= "00000111000000000001011100000100";
wait for Clk_period;
Addr <= "0110010111001";
Trees_din <= "00000000000110000011010010001101";
wait for Clk_period;
Addr <= "0110010111010";
Trees_din <= "00000000011001000011010010001101";
wait for Clk_period;
Addr <= "0110010111011";
Trees_din <= "00000011000000000010011000000100";
wait for Clk_period;
Addr <= "0110010111100";
Trees_din <= "00000000001000010011010010001101";
wait for Clk_period;
Addr <= "0110010111101";
Trees_din <= "00000000010101010011010010001101";
wait for Clk_period;
Addr <= "0110010111110";
Trees_din <= "00000000000000000101010100001000";
wait for Clk_period;
Addr <= "0110010111111";
Trees_din <= "00000000000000000010100100000100";
wait for Clk_period;
Addr <= "0110011000000";
Trees_din <= "00000000000100110011010010001101";
wait for Clk_period;
Addr <= "0110011000001";
Trees_din <= "00000000001000000011010010001101";
wait for Clk_period;
Addr <= "0110011000010";
Trees_din <= "00000101000000000010011000000100";
wait for Clk_period;
Addr <= "0110011000011";
Trees_din <= "00000000000111000011010010001101";
wait for Clk_period;
Addr <= "0110011000100";
Trees_din <= "00000000001110000011010010001101";
wait for Clk_period;
Addr <= "0110011000101";
Trees_din <= "00000111000000000110001000100000";
wait for Clk_period;
Addr <= "0110011000110";
Trees_din <= "00000100000000000001001100010000";
wait for Clk_period;
Addr <= "0110011000111";
Trees_din <= "00000010000000000010100100001000";
wait for Clk_period;
Addr <= "0110011001000";
Trees_din <= "00000101000000000010000100000100";
wait for Clk_period;
Addr <= "0110011001001";
Trees_din <= "00000000011000010011010010001101";
wait for Clk_period;
Addr <= "0110011001010";
Trees_din <= "00000000001010100011010010001101";
wait for Clk_period;
Addr <= "0110011001011";
Trees_din <= "00000100000000000010111100000100";
wait for Clk_period;
Addr <= "0110011001100";
Trees_din <= "00000000000110010011010010001101";
wait for Clk_period;
Addr <= "0110011001101";
Trees_din <= "00000000011000000011010010001101";
wait for Clk_period;
Addr <= "0110011001110";
Trees_din <= "00000111000000000010010100001000";
wait for Clk_period;
Addr <= "0110011001111";
Trees_din <= "00000100000000000100110100000100";
wait for Clk_period;
Addr <= "0110011010000";
Trees_din <= "00000000010111010011010010001101";
wait for Clk_period;
Addr <= "0110011010001";
Trees_din <= "00000000001111000011010010001101";
wait for Clk_period;
Addr <= "0110011010010";
Trees_din <= "00000000000000000000111000000100";
wait for Clk_period;
Addr <= "0110011010011";
Trees_din <= "00000000001100110011010010001101";
wait for Clk_period;
Addr <= "0110011010100";
Trees_din <= "00000000001100010011010010001101";
wait for Clk_period;
Addr <= "0110011010101";
Trees_din <= "00000100000000000010101000010000";
wait for Clk_period;
Addr <= "0110011010110";
Trees_din <= "00000100000000000000110100001000";
wait for Clk_period;
Addr <= "0110011010111";
Trees_din <= "00000001000000000000101100000100";
wait for Clk_period;
Addr <= "0110011011000";
Trees_din <= "00000000000010110011010010001101";
wait for Clk_period;
Addr <= "0110011011001";
Trees_din <= "00000000000111100011010010001101";
wait for Clk_period;
Addr <= "0110011011010";
Trees_din <= "00000010000000000101010000000100";
wait for Clk_period;
Addr <= "0110011011011";
Trees_din <= "00000000001000100011010010001101";
wait for Clk_period;
Addr <= "0110011011100";
Trees_din <= "00000000000101100011010010001101";
wait for Clk_period;
Addr <= "0110011011101";
Trees_din <= "00000000000000000101101000001000";
wait for Clk_period;
Addr <= "0110011011110";
Trees_din <= "00000111000000000101000000000100";
wait for Clk_period;
Addr <= "0110011011111";
Trees_din <= "00000000010111010011010010001101";
wait for Clk_period;
Addr <= "0110011100000";
Trees_din <= "00000000001000100011010010001101";
wait for Clk_period;
Addr <= "0110011100001";
Trees_din <= "00000011000000000101011000000100";
wait for Clk_period;
Addr <= "0110011100010";
Trees_din <= "00000000001010000011010010001101";
wait for Clk_period;
Addr <= "0110011100011";
Trees_din <= "00000000010010010011010010001101";
wait for Clk_period;
Addr <= "0110011100100";
Trees_din <= "00000011000000000001011101000000";
wait for Clk_period;
Addr <= "0110011100101";
Trees_din <= "00000000000000000011101000100000";
wait for Clk_period;
Addr <= "0110011100110";
Trees_din <= "00000010000000000011111100010000";
wait for Clk_period;
Addr <= "0110011100111";
Trees_din <= "00000111000000000011111100001000";
wait for Clk_period;
Addr <= "0110011101000";
Trees_din <= "00000001000000000101111100000100";
wait for Clk_period;
Addr <= "0110011101001";
Trees_din <= "00000000001111000011010010001101";
wait for Clk_period;
Addr <= "0110011101010";
Trees_din <= "00000000010100110011010010001101";
wait for Clk_period;
Addr <= "0110011101011";
Trees_din <= "00000100000000000000010000000100";
wait for Clk_period;
Addr <= "0110011101100";
Trees_din <= "00000000010011110011010010001101";
wait for Clk_period;
Addr <= "0110011101101";
Trees_din <= "00000000001011000011010010001101";
wait for Clk_period;
Addr <= "0110011101110";
Trees_din <= "00000111000000000010100000001000";
wait for Clk_period;
Addr <= "0110011101111";
Trees_din <= "00000110000000000000001000000100";
wait for Clk_period;
Addr <= "0110011110000";
Trees_din <= "00000000001110100011010010001101";
wait for Clk_period;
Addr <= "0110011110001";
Trees_din <= "00000000000011010011010010001101";
wait for Clk_period;
Addr <= "0110011110010";
Trees_din <= "00000110000000000011100100000100";
wait for Clk_period;
Addr <= "0110011110011";
Trees_din <= "00000000000110100011010010001101";
wait for Clk_period;
Addr <= "0110011110100";
Trees_din <= "00000000010001000011010010001101";
wait for Clk_period;
Addr <= "0110011110101";
Trees_din <= "00000110000000000000011100010000";
wait for Clk_period;
Addr <= "0110011110110";
Trees_din <= "00000101000000000101000100001000";
wait for Clk_period;
Addr <= "0110011110111";
Trees_din <= "00000101000000000011100000000100";
wait for Clk_period;
Addr <= "0110011111000";
Trees_din <= "00000000010111000011010010001101";
wait for Clk_period;
Addr <= "0110011111001";
Trees_din <= "00000000000110100011010010001101";
wait for Clk_period;
Addr <= "0110011111010";
Trees_din <= "00000101000000000101001100000100";
wait for Clk_period;
Addr <= "0110011111011";
Trees_din <= "00000000001011010011010010001101";
wait for Clk_period;
Addr <= "0110011111100";
Trees_din <= "00000000000111110011010010001101";
wait for Clk_period;
Addr <= "0110011111101";
Trees_din <= "00000001000000000011111100001000";
wait for Clk_period;
Addr <= "0110011111110";
Trees_din <= "00000111000000000011110000000100";
wait for Clk_period;
Addr <= "0110011111111";
Trees_din <= "00000000000011110011010010001101";
wait for Clk_period;
Addr <= "0110100000000";
Trees_din <= "00000000000011010011010010001101";
wait for Clk_period;
Addr <= "0110100000001";
Trees_din <= "00000010000000000011110100000100";
wait for Clk_period;
Addr <= "0110100000010";
Trees_din <= "00000000001101100011010010001101";
wait for Clk_period;
Addr <= "0110100000011";
Trees_din <= "00000000000101110011010010001101";
wait for Clk_period;
Addr <= "0110100000100";
Trees_din <= "00000110000000000011110000100000";
wait for Clk_period;
Addr <= "0110100000101";
Trees_din <= "00000111000000000110001100010000";
wait for Clk_period;
Addr <= "0110100000110";
Trees_din <= "00000101000000000101100000001000";
wait for Clk_period;
Addr <= "0110100000111";
Trees_din <= "00000001000000000101000100000100";
wait for Clk_period;
Addr <= "0110100001000";
Trees_din <= "00000000011000010011010010001101";
wait for Clk_period;
Addr <= "0110100001001";
Trees_din <= "00000000000000100011010010001101";
wait for Clk_period;
Addr <= "0110100001010";
Trees_din <= "00000100000000000001001100000100";
wait for Clk_period;
Addr <= "0110100001011";
Trees_din <= "00000000001101010011010010001101";
wait for Clk_period;
Addr <= "0110100001100";
Trees_din <= "00000000010001000011010010001101";
wait for Clk_period;
Addr <= "0110100001101";
Trees_din <= "00000011000000000100101000001000";
wait for Clk_period;
Addr <= "0110100001110";
Trees_din <= "00000101000000000000110100000100";
wait for Clk_period;
Addr <= "0110100001111";
Trees_din <= "00000000010100100011010010001101";
wait for Clk_period;
Addr <= "0110100010000";
Trees_din <= "00000000001100110011010010001101";
wait for Clk_period;
Addr <= "0110100010001";
Trees_din <= "00000101000000000101101100000100";
wait for Clk_period;
Addr <= "0110100010010";
Trees_din <= "00000000000111100011010010001101";
wait for Clk_period;
Addr <= "0110100010011";
Trees_din <= "00000000001010000011010010001101";
wait for Clk_period;
Addr <= "0110100010100";
Trees_din <= "00000100000000000101101000010000";
wait for Clk_period;
Addr <= "0110100010101";
Trees_din <= "00000000000000000001110000001000";
wait for Clk_period;
Addr <= "0110100010110";
Trees_din <= "00000010000000000101010000000100";
wait for Clk_period;
Addr <= "0110100010111";
Trees_din <= "00000000001011110011010010001101";
wait for Clk_period;
Addr <= "0110100011000";
Trees_din <= "00000000010010100011010010001101";
wait for Clk_period;
Addr <= "0110100011001";
Trees_din <= "00000010000000000100010100000100";
wait for Clk_period;
Addr <= "0110100011010";
Trees_din <= "00000000010000010011010010001101";
wait for Clk_period;
Addr <= "0110100011011";
Trees_din <= "00000000001000000011010010001101";
wait for Clk_period;
Addr <= "0110100011100";
Trees_din <= "00000111000000000011000100001000";
wait for Clk_period;
Addr <= "0110100011101";
Trees_din <= "00000000000000000001100000000100";
wait for Clk_period;
Addr <= "0110100011110";
Trees_din <= "00000000001111100011010010001101";
wait for Clk_period;
Addr <= "0110100011111";
Trees_din <= "00000000010110000011010010001101";
wait for Clk_period;
Addr <= "0110100100000";
Trees_din <= "00000011000000000101110100000100";
wait for Clk_period;
Addr <= "0110100100001";
Trees_din <= "00000000000101100011010010001101";
wait for Clk_period;
Addr <= "0110100100010";
Trees_din <= "00000000010011100011010010001101";
wait for Clk_period;



----------tree 26-------------------

Addr <= "0110100100011";
Trees_din <= "00000100000000000001110110000000";
wait for Clk_period;
Addr <= "0110100100100";
Trees_din <= "00000001000000000001011001000000";
wait for Clk_period;
Addr <= "0110100100101";
Trees_din <= "00000000000000000010100000100000";
wait for Clk_period;
Addr <= "0110100100110";
Trees_din <= "00000001000000000101001100010000";
wait for Clk_period;
Addr <= "0110100100111";
Trees_din <= "00000000000000000100111000001000";
wait for Clk_period;
Addr <= "0110100101000";
Trees_din <= "00000111000000000101010100000100";
wait for Clk_period;
Addr <= "0110100101001";
Trees_din <= "00000000001110110011011010001001";
wait for Clk_period;
Addr <= "0110100101010";
Trees_din <= "00000000010110110011011010001001";
wait for Clk_period;
Addr <= "0110100101011";
Trees_din <= "00000010000000000010000100000100";
wait for Clk_period;
Addr <= "0110100101100";
Trees_din <= "00000000000101110011011010001001";
wait for Clk_period;
Addr <= "0110100101101";
Trees_din <= "00000000000000110011011010001001";
wait for Clk_period;
Addr <= "0110100101110";
Trees_din <= "00000001000000000101110100001000";
wait for Clk_period;
Addr <= "0110100101111";
Trees_din <= "00000001000000000000111100000100";
wait for Clk_period;
Addr <= "0110100110000";
Trees_din <= "00000000001110000011011010001001";
wait for Clk_period;
Addr <= "0110100110001";
Trees_din <= "00000000001101100011011010001001";
wait for Clk_period;
Addr <= "0110100110010";
Trees_din <= "00000100000000000010110100000100";
wait for Clk_period;
Addr <= "0110100110011";
Trees_din <= "00000000000100100011011010001001";
wait for Clk_period;
Addr <= "0110100110100";
Trees_din <= "00000000011001000011011010001001";
wait for Clk_period;
Addr <= "0110100110101";
Trees_din <= "00000100000000000010100000010000";
wait for Clk_period;
Addr <= "0110100110110";
Trees_din <= "00000010000000000010110100001000";
wait for Clk_period;
Addr <= "0110100110111";
Trees_din <= "00000101000000000001011100000100";
wait for Clk_period;
Addr <= "0110100111000";
Trees_din <= "00000000001101010011011010001001";
wait for Clk_period;
Addr <= "0110100111001";
Trees_din <= "00000000001001110011011010001001";
wait for Clk_period;
Addr <= "0110100111010";
Trees_din <= "00000011000000000100100100000100";
wait for Clk_period;
Addr <= "0110100111011";
Trees_din <= "00000000000001110011011010001001";
wait for Clk_period;
Addr <= "0110100111100";
Trees_din <= "00000000000101000011011010001001";
wait for Clk_period;
Addr <= "0110100111101";
Trees_din <= "00000100000000000100011000001000";
wait for Clk_period;
Addr <= "0110100111110";
Trees_din <= "00000100000000000010011000000100";
wait for Clk_period;
Addr <= "0110100111111";
Trees_din <= "00000000000010100011011010001001";
wait for Clk_period;
Addr <= "0110101000000";
Trees_din <= "00000000000101010011011010001001";
wait for Clk_period;
Addr <= "0110101000001";
Trees_din <= "00000000000000000101001100000100";
wait for Clk_period;
Addr <= "0110101000010";
Trees_din <= "00000000000000110011011010001001";
wait for Clk_period;
Addr <= "0110101000011";
Trees_din <= "00000000010100000011011010001001";
wait for Clk_period;
Addr <= "0110101000100";
Trees_din <= "00000010000000000000111100100000";
wait for Clk_period;
Addr <= "0110101000101";
Trees_din <= "00000111000000000011011100010000";
wait for Clk_period;
Addr <= "0110101000110";
Trees_din <= "00000010000000000000010000001000";
wait for Clk_period;
Addr <= "0110101000111";
Trees_din <= "00000110000000000010100000000100";
wait for Clk_period;
Addr <= "0110101001000";
Trees_din <= "00000000000101100011011010001001";
wait for Clk_period;
Addr <= "0110101001001";
Trees_din <= "00000000001110000011011010001001";
wait for Clk_period;
Addr <= "0110101001010";
Trees_din <= "00000001000000000100110000000100";
wait for Clk_period;
Addr <= "0110101001011";
Trees_din <= "00000000000000110011011010001001";
wait for Clk_period;
Addr <= "0110101001100";
Trees_din <= "00000000011000100011011010001001";
wait for Clk_period;
Addr <= "0110101001101";
Trees_din <= "00000001000000000101101100001000";
wait for Clk_period;
Addr <= "0110101001110";
Trees_din <= "00000011000000000010011100000100";
wait for Clk_period;
Addr <= "0110101001111";
Trees_din <= "00000000011000100011011010001001";
wait for Clk_period;
Addr <= "0110101010000";
Trees_din <= "00000000001001110011011010001001";
wait for Clk_period;
Addr <= "0110101010001";
Trees_din <= "00000110000000000101101000000100";
wait for Clk_period;
Addr <= "0110101010010";
Trees_din <= "00000000010111110011011010001001";
wait for Clk_period;
Addr <= "0110101010011";
Trees_din <= "00000000001100100011011010001001";
wait for Clk_period;
Addr <= "0110101010100";
Trees_din <= "00000001000000000001000100010000";
wait for Clk_period;
Addr <= "0110101010101";
Trees_din <= "00000011000000000101001000001000";
wait for Clk_period;
Addr <= "0110101010110";
Trees_din <= "00000101000000000011101000000100";
wait for Clk_period;
Addr <= "0110101010111";
Trees_din <= "00000000000000010011011010001001";
wait for Clk_period;
Addr <= "0110101011000";
Trees_din <= "00000000001100000011011010001001";
wait for Clk_period;
Addr <= "0110101011001";
Trees_din <= "00000000000000000100100000000100";
wait for Clk_period;
Addr <= "0110101011010";
Trees_din <= "00000000000100000011011010001001";
wait for Clk_period;
Addr <= "0110101011011";
Trees_din <= "00000000001011110011011010001001";
wait for Clk_period;
Addr <= "0110101011100";
Trees_din <= "00000011000000000010010100001000";
wait for Clk_period;
Addr <= "0110101011101";
Trees_din <= "00000000000000000101111100000100";
wait for Clk_period;
Addr <= "0110101011110";
Trees_din <= "00000000010000000011011010001001";
wait for Clk_period;
Addr <= "0110101011111";
Trees_din <= "00000000001101000011011010001001";
wait for Clk_period;
Addr <= "0110101100000";
Trees_din <= "00000100000000000101111000000100";
wait for Clk_period;
Addr <= "0110101100001";
Trees_din <= "00000000000001010011011010001001";
wait for Clk_period;
Addr <= "0110101100010";
Trees_din <= "00000000001100110011011010001001";
wait for Clk_period;
Addr <= "0110101100011";
Trees_din <= "00000000000000000101001101000000";
wait for Clk_period;
Addr <= "0110101100100";
Trees_din <= "00000110000000000100100000100000";
wait for Clk_period;
Addr <= "0110101100101";
Trees_din <= "00000111000000000100000000010000";
wait for Clk_period;
Addr <= "0110101100110";
Trees_din <= "00000011000000000000010100001000";
wait for Clk_period;
Addr <= "0110101100111";
Trees_din <= "00000100000000000000100000000100";
wait for Clk_period;
Addr <= "0110101101000";
Trees_din <= "00000000000000000011011010001001";
wait for Clk_period;
Addr <= "0110101101001";
Trees_din <= "00000000011000100011011010001001";
wait for Clk_period;
Addr <= "0110101101010";
Trees_din <= "00000101000000000100000000000100";
wait for Clk_period;
Addr <= "0110101101011";
Trees_din <= "00000000000110110011011010001001";
wait for Clk_period;
Addr <= "0110101101100";
Trees_din <= "00000000000111100011011010001001";
wait for Clk_period;
Addr <= "0110101101101";
Trees_din <= "00000110000000000000000000001000";
wait for Clk_period;
Addr <= "0110101101110";
Trees_din <= "00000100000000000000110000000100";
wait for Clk_period;
Addr <= "0110101101111";
Trees_din <= "00000000001100010011011010001001";
wait for Clk_period;
Addr <= "0110101110000";
Trees_din <= "00000000000100100011011010001001";
wait for Clk_period;
Addr <= "0110101110001";
Trees_din <= "00000000000000000011000000000100";
wait for Clk_period;
Addr <= "0110101110010";
Trees_din <= "00000000001011010011011010001001";
wait for Clk_period;
Addr <= "0110101110011";
Trees_din <= "00000000000000110011011010001001";
wait for Clk_period;
Addr <= "0110101110100";
Trees_din <= "00000111000000000011100100010000";
wait for Clk_period;
Addr <= "0110101110101";
Trees_din <= "00000100000000000001110100001000";
wait for Clk_period;
Addr <= "0110101110110";
Trees_din <= "00000111000000000000000000000100";
wait for Clk_period;
Addr <= "0110101110111";
Trees_din <= "00000000000111000011011010001001";
wait for Clk_period;
Addr <= "0110101111000";
Trees_din <= "00000000000111100011011010001001";
wait for Clk_period;
Addr <= "0110101111001";
Trees_din <= "00000000000000000101001000000100";
wait for Clk_period;
Addr <= "0110101111010";
Trees_din <= "00000000010101000011011010001001";
wait for Clk_period;
Addr <= "0110101111011";
Trees_din <= "00000000000111010011011010001001";
wait for Clk_period;
Addr <= "0110101111100";
Trees_din <= "00000110000000000100011000001000";
wait for Clk_period;
Addr <= "0110101111101";
Trees_din <= "00000011000000000010011100000100";
wait for Clk_period;
Addr <= "0110101111110";
Trees_din <= "00000000000011000011011010001001";
wait for Clk_period;
Addr <= "0110101111111";
Trees_din <= "00000000001111000011011010001001";
wait for Clk_period;
Addr <= "0110110000000";
Trees_din <= "00000011000000000100111000000100";
wait for Clk_period;
Addr <= "0110110000001";
Trees_din <= "00000000001111110011011010001001";
wait for Clk_period;
Addr <= "0110110000010";
Trees_din <= "00000000000111000011011010001001";
wait for Clk_period;
Addr <= "0110110000011";
Trees_din <= "00000100000000000101001100100000";
wait for Clk_period;
Addr <= "0110110000100";
Trees_din <= "00000010000000000001111100010000";
wait for Clk_period;
Addr <= "0110110000101";
Trees_din <= "00000110000000000100011100001000";
wait for Clk_period;
Addr <= "0110110000110";
Trees_din <= "00000101000000000010111000000100";
wait for Clk_period;
Addr <= "0110110000111";
Trees_din <= "00000000001110110011011010001001";
wait for Clk_period;
Addr <= "0110110001000";
Trees_din <= "00000000000110100011011010001001";
wait for Clk_period;
Addr <= "0110110001001";
Trees_din <= "00000101000000000010110100000100";
wait for Clk_period;
Addr <= "0110110001010";
Trees_din <= "00000000010001110011011010001001";
wait for Clk_period;
Addr <= "0110110001011";
Trees_din <= "00000000001111010011011010001001";
wait for Clk_period;
Addr <= "0110110001100";
Trees_din <= "00000101000000000101111000001000";
wait for Clk_period;
Addr <= "0110110001101";
Trees_din <= "00000110000000000010010100000100";
wait for Clk_period;
Addr <= "0110110001110";
Trees_din <= "00000000001110110011011010001001";
wait for Clk_period;
Addr <= "0110110001111";
Trees_din <= "00000000010001100011011010001001";
wait for Clk_period;
Addr <= "0110110010000";
Trees_din <= "00000111000000000011111100000100";
wait for Clk_period;
Addr <= "0110110010001";
Trees_din <= "00000000001101010011011010001001";
wait for Clk_period;
Addr <= "0110110010010";
Trees_din <= "00000000001111000011011010001001";
wait for Clk_period;
Addr <= "0110110010011";
Trees_din <= "00000111000000000010001100010000";
wait for Clk_period;
Addr <= "0110110010100";
Trees_din <= "00000101000000000011101100001000";
wait for Clk_period;
Addr <= "0110110010101";
Trees_din <= "00000101000000000110000100000100";
wait for Clk_period;
Addr <= "0110110010110";
Trees_din <= "00000000001100110011011010001001";
wait for Clk_period;
Addr <= "0110110010111";
Trees_din <= "00000000001011110011011010001001";
wait for Clk_period;
Addr <= "0110110011000";
Trees_din <= "00000000000000000100111000000100";
wait for Clk_period;
Addr <= "0110110011001";
Trees_din <= "00000000000001000011011010001001";
wait for Clk_period;
Addr <= "0110110011010";
Trees_din <= "00000000001100100011011010001001";
wait for Clk_period;
Addr <= "0110110011011";
Trees_din <= "00000010000000000011001000001000";
wait for Clk_period;
Addr <= "0110110011100";
Trees_din <= "00000001000000000101011100000100";
wait for Clk_period;
Addr <= "0110110011101";
Trees_din <= "00000000011000010011011010001001";
wait for Clk_period;
Addr <= "0110110011110";
Trees_din <= "00000000001100010011011010001001";
wait for Clk_period;
Addr <= "0110110011111";
Trees_din <= "00000110000000000010001000000100";
wait for Clk_period;
Addr <= "0110110100000";
Trees_din <= "00000000001010010011011010001001";
wait for Clk_period;
Addr <= "0110110100001";
Trees_din <= "00000000000111000011011010001001";
wait for Clk_period;



----------tree 27-------------------

Addr <= "0110110100010";
Trees_din <= "00000001000000000010111010000000";
wait for Clk_period;
Addr <= "0110110100011";
Trees_din <= "00000001000000000000000101000000";
wait for Clk_period;
Addr <= "0110110100100";
Trees_din <= "00000110000000000010101100100000";
wait for Clk_period;
Addr <= "0110110100101";
Trees_din <= "00000110000000000000110000010000";
wait for Clk_period;
Addr <= "0110110100110";
Trees_din <= "00000110000000000101110000001000";
wait for Clk_period;
Addr <= "0110110100111";
Trees_din <= "00000110000000000110000100000100";
wait for Clk_period;
Addr <= "0110110101000";
Trees_din <= "00000000010011110011100010000101";
wait for Clk_period;
Addr <= "0110110101001";
Trees_din <= "00000000000010000011100010000101";
wait for Clk_period;
Addr <= "0110110101010";
Trees_din <= "00000001000000000001000100000100";
wait for Clk_period;
Addr <= "0110110101011";
Trees_din <= "00000000001011110011100010000101";
wait for Clk_period;
Addr <= "0110110101100";
Trees_din <= "00000000000110100011100010000101";
wait for Clk_period;
Addr <= "0110110101101";
Trees_din <= "00000010000000000000011000001000";
wait for Clk_period;
Addr <= "0110110101110";
Trees_din <= "00000100000000000000011100000100";
wait for Clk_period;
Addr <= "0110110101111";
Trees_din <= "00000000000010000011100010000101";
wait for Clk_period;
Addr <= "0110110110000";
Trees_din <= "00000000001111100011100010000101";
wait for Clk_period;
Addr <= "0110110110001";
Trees_din <= "00000100000000000010111000000100";
wait for Clk_period;
Addr <= "0110110110010";
Trees_din <= "00000000001010100011100010000101";
wait for Clk_period;
Addr <= "0110110110011";
Trees_din <= "00000000000010110011100010000101";
wait for Clk_period;
Addr <= "0110110110100";
Trees_din <= "00000011000000000010010100010000";
wait for Clk_period;
Addr <= "0110110110101";
Trees_din <= "00000100000000000100010000001000";
wait for Clk_period;
Addr <= "0110110110110";
Trees_din <= "00000010000000000001111000000100";
wait for Clk_period;
Addr <= "0110110110111";
Trees_din <= "00000000001010100011100010000101";
wait for Clk_period;
Addr <= "0110110111000";
Trees_din <= "00000000000110100011100010000101";
wait for Clk_period;
Addr <= "0110110111001";
Trees_din <= "00000011000000000010010100000100";
wait for Clk_period;
Addr <= "0110110111010";
Trees_din <= "00000000000001010011100010000101";
wait for Clk_period;
Addr <= "0110110111011";
Trees_din <= "00000000000110000011100010000101";
wait for Clk_period;
Addr <= "0110110111100";
Trees_din <= "00000110000000000101111000001000";
wait for Clk_period;
Addr <= "0110110111101";
Trees_din <= "00000110000000000000110100000100";
wait for Clk_period;
Addr <= "0110110111110";
Trees_din <= "00000000001100110011100010000101";
wait for Clk_period;
Addr <= "0110110111111";
Trees_din <= "00000000001011000011100010000101";
wait for Clk_period;
Addr <= "0110111000000";
Trees_din <= "00000101000000000011101100000100";
wait for Clk_period;
Addr <= "0110111000001";
Trees_din <= "00000000000111110011100010000101";
wait for Clk_period;
Addr <= "0110111000010";
Trees_din <= "00000000001001010011100010000101";
wait for Clk_period;
Addr <= "0110111000011";
Trees_din <= "00000001000000000011010000100000";
wait for Clk_period;
Addr <= "0110111000100";
Trees_din <= "00000000000000000010001100010000";
wait for Clk_period;
Addr <= "0110111000101";
Trees_din <= "00000010000000000001001100001000";
wait for Clk_period;
Addr <= "0110111000110";
Trees_din <= "00000100000000000100100000000100";
wait for Clk_period;
Addr <= "0110111000111";
Trees_din <= "00000000010000000011100010000101";
wait for Clk_period;
Addr <= "0110111001000";
Trees_din <= "00000000000110010011100010000101";
wait for Clk_period;
Addr <= "0110111001001";
Trees_din <= "00000001000000000101011000000100";
wait for Clk_period;
Addr <= "0110111001010";
Trees_din <= "00000000010110110011100010000101";
wait for Clk_period;
Addr <= "0110111001011";
Trees_din <= "00000000010110100011100010000101";
wait for Clk_period;
Addr <= "0110111001100";
Trees_din <= "00000011000000000011000000001000";
wait for Clk_period;
Addr <= "0110111001101";
Trees_din <= "00000000000000000101101100000100";
wait for Clk_period;
Addr <= "0110111001110";
Trees_din <= "00000000000110010011100010000101";
wait for Clk_period;
Addr <= "0110111001111";
Trees_din <= "00000000000110000011100010000101";
wait for Clk_period;
Addr <= "0110111010000";
Trees_din <= "00000111000000000101001000000100";
wait for Clk_period;
Addr <= "0110111010001";
Trees_din <= "00000000011000110011100010000101";
wait for Clk_period;
Addr <= "0110111010010";
Trees_din <= "00000000001111000011100010000101";
wait for Clk_period;
Addr <= "0110111010011";
Trees_din <= "00000100000000000001011100010000";
wait for Clk_period;
Addr <= "0110111010100";
Trees_din <= "00000011000000000101000100001000";
wait for Clk_period;
Addr <= "0110111010101";
Trees_din <= "00000110000000000101011100000100";
wait for Clk_period;
Addr <= "0110111010110";
Trees_din <= "00000000000011100011100010000101";
wait for Clk_period;
Addr <= "0110111010111";
Trees_din <= "00000000001100110011100010000101";
wait for Clk_period;
Addr <= "0110111011000";
Trees_din <= "00000100000000000010101100000100";
wait for Clk_period;
Addr <= "0110111011001";
Trees_din <= "00000000000011000011100010000101";
wait for Clk_period;
Addr <= "0110111011010";
Trees_din <= "00000000001110100011100010000101";
wait for Clk_period;
Addr <= "0110111011011";
Trees_din <= "00000101000000000001000000001000";
wait for Clk_period;
Addr <= "0110111011100";
Trees_din <= "00000110000000000010011000000100";
wait for Clk_period;
Addr <= "0110111011101";
Trees_din <= "00000000001101100011100010000101";
wait for Clk_period;
Addr <= "0110111011110";
Trees_din <= "00000000001110010011100010000101";
wait for Clk_period;
Addr <= "0110111011111";
Trees_din <= "00000011000000000110001100000100";
wait for Clk_period;
Addr <= "0110111100000";
Trees_din <= "00000000001100100011100010000101";
wait for Clk_period;
Addr <= "0110111100001";
Trees_din <= "00000000001111010011100010000101";
wait for Clk_period;
Addr <= "0110111100010";
Trees_din <= "00000010000000000001011101000000";
wait for Clk_period;
Addr <= "0110111100011";
Trees_din <= "00000011000000000001001100100000";
wait for Clk_period;
Addr <= "0110111100100";
Trees_din <= "00000111000000000010010000010000";
wait for Clk_period;
Addr <= "0110111100101";
Trees_din <= "00000011000000000110001000001000";
wait for Clk_period;
Addr <= "0110111100110";
Trees_din <= "00000100000000000000100000000100";
wait for Clk_period;
Addr <= "0110111100111";
Trees_din <= "00000000001011000011100010000101";
wait for Clk_period;
Addr <= "0110111101000";
Trees_din <= "00000000010110100011100010000101";
wait for Clk_period;
Addr <= "0110111101001";
Trees_din <= "00000111000000000101011000000100";
wait for Clk_period;
Addr <= "0110111101010";
Trees_din <= "00000000010001010011100010000101";
wait for Clk_period;
Addr <= "0110111101011";
Trees_din <= "00000000010101010011100010000101";
wait for Clk_period;
Addr <= "0110111101100";
Trees_din <= "00000010000000000110000100001000";
wait for Clk_period;
Addr <= "0110111101101";
Trees_din <= "00000001000000000101000100000100";
wait for Clk_period;
Addr <= "0110111101110";
Trees_din <= "00000000010000000011100010000101";
wait for Clk_period;
Addr <= "0110111101111";
Trees_din <= "00000000001101010011100010000101";
wait for Clk_period;
Addr <= "0110111110000";
Trees_din <= "00000011000000000010000000000100";
wait for Clk_period;
Addr <= "0110111110001";
Trees_din <= "00000000000000000011100010000101";
wait for Clk_period;
Addr <= "0110111110010";
Trees_din <= "00000000010110010011100010000101";
wait for Clk_period;
Addr <= "0110111110011";
Trees_din <= "00000111000000000011001100010000";
wait for Clk_period;
Addr <= "0110111110100";
Trees_din <= "00000000000000000100110100001000";
wait for Clk_period;
Addr <= "0110111110101";
Trees_din <= "00000111000000000000100000000100";
wait for Clk_period;
Addr <= "0110111110110";
Trees_din <= "00000000000101100011100010000101";
wait for Clk_period;
Addr <= "0110111110111";
Trees_din <= "00000000000101000011100010000101";
wait for Clk_period;
Addr <= "0110111111000";
Trees_din <= "00000000000000000100100000000100";
wait for Clk_period;
Addr <= "0110111111001";
Trees_din <= "00000000000110010011100010000101";
wait for Clk_period;
Addr <= "0110111111010";
Trees_din <= "00000000000011110011100010000101";
wait for Clk_period;
Addr <= "0110111111011";
Trees_din <= "00000111000000000011011100001000";
wait for Clk_period;
Addr <= "0110111111100";
Trees_din <= "00000011000000000000001000000100";
wait for Clk_period;
Addr <= "0110111111101";
Trees_din <= "00000000000110100011100010000101";
wait for Clk_period;
Addr <= "0110111111110";
Trees_din <= "00000000000100010011100010000101";
wait for Clk_period;
Addr <= "0110111111111";
Trees_din <= "00000101000000000100001000000100";
wait for Clk_period;
Addr <= "0111000000000";
Trees_din <= "00000000010010110011100010000101";
wait for Clk_period;
Addr <= "0111000000001";
Trees_din <= "00000000010000110011100010000101";
wait for Clk_period;
Addr <= "0111000000010";
Trees_din <= "00000011000000000101101000100000";
wait for Clk_period;
Addr <= "0111000000011";
Trees_din <= "00000100000000000000011100010000";
wait for Clk_period;
Addr <= "0111000000100";
Trees_din <= "00000010000000000101101100001000";
wait for Clk_period;
Addr <= "0111000000101";
Trees_din <= "00000011000000000100001000000100";
wait for Clk_period;
Addr <= "0111000000110";
Trees_din <= "00000000010001000011100010000101";
wait for Clk_period;
Addr <= "0111000000111";
Trees_din <= "00000000000011110011100010000101";
wait for Clk_period;
Addr <= "0111000001000";
Trees_din <= "00000000000000000101000100000100";
wait for Clk_period;
Addr <= "0111000001001";
Trees_din <= "00000000000101110011100010000101";
wait for Clk_period;
Addr <= "0111000001010";
Trees_din <= "00000000001101010011100010000101";
wait for Clk_period;
Addr <= "0111000001011";
Trees_din <= "00000110000000000100000000001000";
wait for Clk_period;
Addr <= "0111000001100";
Trees_din <= "00000001000000000010100000000100";
wait for Clk_period;
Addr <= "0111000001101";
Trees_din <= "00000000000000010011100010000101";
wait for Clk_period;
Addr <= "0111000001110";
Trees_din <= "00000000010110110011100010000101";
wait for Clk_period;
Addr <= "0111000001111";
Trees_din <= "00000110000000000001000000000100";
wait for Clk_period;
Addr <= "0111000010000";
Trees_din <= "00000000001010100011100010000101";
wait for Clk_period;
Addr <= "0111000010001";
Trees_din <= "00000000000111100011100010000101";
wait for Clk_period;
Addr <= "0111000010010";
Trees_din <= "00000110000000000011010100010000";
wait for Clk_period;
Addr <= "0111000010011";
Trees_din <= "00000011000000000001101000001000";
wait for Clk_period;
Addr <= "0111000010100";
Trees_din <= "00000001000000000010001100000100";
wait for Clk_period;
Addr <= "0111000010101";
Trees_din <= "00000000011000010011100010000101";
wait for Clk_period;
Addr <= "0111000010110";
Trees_din <= "00000000010111110011100010000101";
wait for Clk_period;
Addr <= "0111000010111";
Trees_din <= "00000011000000000101011000000100";
wait for Clk_period;
Addr <= "0111000011000";
Trees_din <= "00000000000101010011100010000101";
wait for Clk_period;
Addr <= "0111000011001";
Trees_din <= "00000000000110100011100010000101";
wait for Clk_period;
Addr <= "0111000011010";
Trees_din <= "00000111000000000110001100001000";
wait for Clk_period;
Addr <= "0111000011011";
Trees_din <= "00000011000000000110000100000100";
wait for Clk_period;
Addr <= "0111000011100";
Trees_din <= "00000000001100110011100010000101";
wait for Clk_period;
Addr <= "0111000011101";
Trees_din <= "00000000001101100011100010000101";
wait for Clk_period;
Addr <= "0111000011110";
Trees_din <= "00000000000000000010001000000100";
wait for Clk_period;
Addr <= "0111000011111";
Trees_din <= "00000000000101100011100010000101";
wait for Clk_period;
Addr <= "0111000100000";
Trees_din <= "00000000000000110011100010000101";
wait for Clk_period;



----------tree 28-------------------

Addr <= "0111000100001";
Trees_din <= "00000011000000000101001110000000";
wait for Clk_period;
Addr <= "0111000100010";
Trees_din <= "00000100000000000100001001000000";
wait for Clk_period;
Addr <= "0111000100011";
Trees_din <= "00000000000000000000001100100000";
wait for Clk_period;
Addr <= "0111000100100";
Trees_din <= "00000111000000000010001000010000";
wait for Clk_period;
Addr <= "0111000100101";
Trees_din <= "00000111000000000000010000001000";
wait for Clk_period;
Addr <= "0111000100110";
Trees_din <= "00000101000000000100000100000100";
wait for Clk_period;
Addr <= "0111000100111";
Trees_din <= "00000000011000010011101010000001";
wait for Clk_period;
Addr <= "0111000101000";
Trees_din <= "00000000000011110011101010000001";
wait for Clk_period;
Addr <= "0111000101001";
Trees_din <= "00000100000000000011110000000100";
wait for Clk_period;
Addr <= "0111000101010";
Trees_din <= "00000000010110100011101010000001";
wait for Clk_period;
Addr <= "0111000101011";
Trees_din <= "00000000000011110011101010000001";
wait for Clk_period;
Addr <= "0111000101100";
Trees_din <= "00000100000000000011011100001000";
wait for Clk_period;
Addr <= "0111000101101";
Trees_din <= "00000101000000000011111000000100";
wait for Clk_period;
Addr <= "0111000101110";
Trees_din <= "00000000001110010011101010000001";
wait for Clk_period;
Addr <= "0111000101111";
Trees_din <= "00000000010001000011101010000001";
wait for Clk_period;
Addr <= "0111000110000";
Trees_din <= "00000101000000000000011000000100";
wait for Clk_period;
Addr <= "0111000110001";
Trees_din <= "00000000000000010011101010000001";
wait for Clk_period;
Addr <= "0111000110010";
Trees_din <= "00000000001101110011101010000001";
wait for Clk_period;
Addr <= "0111000110011";
Trees_din <= "00000101000000000011100000010000";
wait for Clk_period;
Addr <= "0111000110100";
Trees_din <= "00000001000000000000101100001000";
wait for Clk_period;
Addr <= "0111000110101";
Trees_din <= "00000010000000000101111100000100";
wait for Clk_period;
Addr <= "0111000110110";
Trees_din <= "00000000010100110011101010000001";
wait for Clk_period;
Addr <= "0111000110111";
Trees_din <= "00000000001010100011101010000001";
wait for Clk_period;
Addr <= "0111000111000";
Trees_din <= "00000000000000000110010000000100";
wait for Clk_period;
Addr <= "0111000111001";
Trees_din <= "00000000001110110011101010000001";
wait for Clk_period;
Addr <= "0111000111010";
Trees_din <= "00000000001000100011101010000001";
wait for Clk_period;
Addr <= "0111000111011";
Trees_din <= "00000010000000000100010100001000";
wait for Clk_period;
Addr <= "0111000111100";
Trees_din <= "00000000000000000101101100000100";
wait for Clk_period;
Addr <= "0111000111101";
Trees_din <= "00000000011000110011101010000001";
wait for Clk_period;
Addr <= "0111000111110";
Trees_din <= "00000000010010000011101010000001";
wait for Clk_period;
Addr <= "0111000111111";
Trees_din <= "00000101000000000010001000000100";
wait for Clk_period;
Addr <= "0111001000000";
Trees_din <= "00000000001000000011101010000001";
wait for Clk_period;
Addr <= "0111001000001";
Trees_din <= "00000000000001010011101010000001";
wait for Clk_period;
Addr <= "0111001000010";
Trees_din <= "00000000000000000100001000100000";
wait for Clk_period;
Addr <= "0111001000011";
Trees_din <= "00000101000000000100111000010000";
wait for Clk_period;
Addr <= "0111001000100";
Trees_din <= "00000100000000000000101000001000";
wait for Clk_period;
Addr <= "0111001000101";
Trees_din <= "00000111000000000010001000000100";
wait for Clk_period;
Addr <= "0111001000110";
Trees_din <= "00000000000001010011101010000001";
wait for Clk_period;
Addr <= "0111001000111";
Trees_din <= "00000000000011010011101010000001";
wait for Clk_period;
Addr <= "0111001001000";
Trees_din <= "00000011000000000101010000000100";
wait for Clk_period;
Addr <= "0111001001001";
Trees_din <= "00000000001010100011101010000001";
wait for Clk_period;
Addr <= "0111001001010";
Trees_din <= "00000000000110010011101010000001";
wait for Clk_period;
Addr <= "0111001001011";
Trees_din <= "00000001000000000011001100001000";
wait for Clk_period;
Addr <= "0111001001100";
Trees_din <= "00000011000000000101000000000100";
wait for Clk_period;
Addr <= "0111001001101";
Trees_din <= "00000000000000110011101010000001";
wait for Clk_period;
Addr <= "0111001001110";
Trees_din <= "00000000010001100011101010000001";
wait for Clk_period;
Addr <= "0111001001111";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "0111001010000";
Trees_din <= "00000000001000010011101010000001";
wait for Clk_period;
Addr <= "0111001010001";
Trees_din <= "00000000001001000011101010000001";
wait for Clk_period;
Addr <= "0111001010010";
Trees_din <= "00000110000000000001101000010000";
wait for Clk_period;
Addr <= "0111001010011";
Trees_din <= "00000110000000000011110100001000";
wait for Clk_period;
Addr <= "0111001010100";
Trees_din <= "00000101000000000101110100000100";
wait for Clk_period;
Addr <= "0111001010101";
Trees_din <= "00000000000011110011101010000001";
wait for Clk_period;
Addr <= "0111001010110";
Trees_din <= "00000000001110010011101010000001";
wait for Clk_period;
Addr <= "0111001010111";
Trees_din <= "00000001000000000011001100000100";
wait for Clk_period;
Addr <= "0111001011000";
Trees_din <= "00000000001100110011101010000001";
wait for Clk_period;
Addr <= "0111001011001";
Trees_din <= "00000000010000100011101010000001";
wait for Clk_period;
Addr <= "0111001011010";
Trees_din <= "00000001000000000000100100001000";
wait for Clk_period;
Addr <= "0111001011011";
Trees_din <= "00000101000000000011100100000100";
wait for Clk_period;
Addr <= "0111001011100";
Trees_din <= "00000000010111010011101010000001";
wait for Clk_period;
Addr <= "0111001011101";
Trees_din <= "00000000001100010011101010000001";
wait for Clk_period;
Addr <= "0111001011110";
Trees_din <= "00000101000000000011011100000100";
wait for Clk_period;
Addr <= "0111001011111";
Trees_din <= "00000000000101100011101010000001";
wait for Clk_period;
Addr <= "0111001100000";
Trees_din <= "00000000010111100011101010000001";
wait for Clk_period;
Addr <= "0111001100001";
Trees_din <= "00000011000000000000101101000000";
wait for Clk_period;
Addr <= "0111001100010";
Trees_din <= "00000110000000000000001100100000";
wait for Clk_period;
Addr <= "0111001100011";
Trees_din <= "00000000000000000000011100010000";
wait for Clk_period;
Addr <= "0111001100100";
Trees_din <= "00000010000000000011001000001000";
wait for Clk_period;
Addr <= "0111001100101";
Trees_din <= "00000010000000000001011000000100";
wait for Clk_period;
Addr <= "0111001100110";
Trees_din <= "00000000001010110011101010000001";
wait for Clk_period;
Addr <= "0111001100111";
Trees_din <= "00000000010011000011101010000001";
wait for Clk_period;
Addr <= "0111001101000";
Trees_din <= "00000110000000000101000000000100";
wait for Clk_period;
Addr <= "0111001101001";
Trees_din <= "00000000001110000011101010000001";
wait for Clk_period;
Addr <= "0111001101010";
Trees_din <= "00000000000001010011101010000001";
wait for Clk_period;
Addr <= "0111001101011";
Trees_din <= "00000101000000000001111100001000";
wait for Clk_period;
Addr <= "0111001101100";
Trees_din <= "00000100000000000010101100000100";
wait for Clk_period;
Addr <= "0111001101101";
Trees_din <= "00000000010000100011101010000001";
wait for Clk_period;
Addr <= "0111001101110";
Trees_din <= "00000000001101110011101010000001";
wait for Clk_period;
Addr <= "0111001101111";
Trees_din <= "00000110000000000110001000000100";
wait for Clk_period;
Addr <= "0111001110000";
Trees_din <= "00000000000101010011101010000001";
wait for Clk_period;
Addr <= "0111001110001";
Trees_din <= "00000000001011110011101010000001";
wait for Clk_period;
Addr <= "0111001110010";
Trees_din <= "00000100000000000011001100010000";
wait for Clk_period;
Addr <= "0111001110011";
Trees_din <= "00000100000000000101100100001000";
wait for Clk_period;
Addr <= "0111001110100";
Trees_din <= "00000001000000000101010100000100";
wait for Clk_period;
Addr <= "0111001110101";
Trees_din <= "00000000001010110011101010000001";
wait for Clk_period;
Addr <= "0111001110110";
Trees_din <= "00000000010000100011101010000001";
wait for Clk_period;
Addr <= "0111001110111";
Trees_din <= "00000001000000000101000100000100";
wait for Clk_period;
Addr <= "0111001111000";
Trees_din <= "00000000001000010011101010000001";
wait for Clk_period;
Addr <= "0111001111001";
Trees_din <= "00000000010101000011101010000001";
wait for Clk_period;
Addr <= "0111001111010";
Trees_din <= "00000111000000000101010100001000";
wait for Clk_period;
Addr <= "0111001111011";
Trees_din <= "00000111000000000000110000000100";
wait for Clk_period;
Addr <= "0111001111100";
Trees_din <= "00000000001111100011101010000001";
wait for Clk_period;
Addr <= "0111001111101";
Trees_din <= "00000000001011100011101010000001";
wait for Clk_period;
Addr <= "0111001111110";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "0111001111111";
Trees_din <= "00000000000011010011101010000001";
wait for Clk_period;
Addr <= "0111010000000";
Trees_din <= "00000000000100010011101010000001";
wait for Clk_period;
Addr <= "0111010000001";
Trees_din <= "00000010000000000011000100100000";
wait for Clk_period;
Addr <= "0111010000010";
Trees_din <= "00000101000000000100011100010000";
wait for Clk_period;
Addr <= "0111010000011";
Trees_din <= "00000001000000000001101000001000";
wait for Clk_period;
Addr <= "0111010000100";
Trees_din <= "00000110000000000001101000000100";
wait for Clk_period;
Addr <= "0111010000101";
Trees_din <= "00000000010111100011101010000001";
wait for Clk_period;
Addr <= "0111010000110";
Trees_din <= "00000000010100110011101010000001";
wait for Clk_period;
Addr <= "0111010000111";
Trees_din <= "00000001000000000000000100000100";
wait for Clk_period;
Addr <= "0111010001000";
Trees_din <= "00000000010111100011101010000001";
wait for Clk_period;
Addr <= "0111010001001";
Trees_din <= "00000000001111000011101010000001";
wait for Clk_period;
Addr <= "0111010001010";
Trees_din <= "00000111000000000101011000001000";
wait for Clk_period;
Addr <= "0111010001011";
Trees_din <= "00000000000000000001000000000100";
wait for Clk_period;
Addr <= "0111010001100";
Trees_din <= "00000000001001000011101010000001";
wait for Clk_period;
Addr <= "0111010001101";
Trees_din <= "00000000000011010011101010000001";
wait for Clk_period;
Addr <= "0111010001110";
Trees_din <= "00000000000000000110001000000100";
wait for Clk_period;
Addr <= "0111010001111";
Trees_din <= "00000000001001010011101010000001";
wait for Clk_period;
Addr <= "0111010010000";
Trees_din <= "00000000001000010011101010000001";
wait for Clk_period;
Addr <= "0111010010001";
Trees_din <= "00000101000000000101100100010000";
wait for Clk_period;
Addr <= "0111010010010";
Trees_din <= "00000101000000000011101100001000";
wait for Clk_period;
Addr <= "0111010010011";
Trees_din <= "00000101000000000000011000000100";
wait for Clk_period;
Addr <= "0111010010100";
Trees_din <= "00000000000001000011101010000001";
wait for Clk_period;
Addr <= "0111010010101";
Trees_din <= "00000000000111110011101010000001";
wait for Clk_period;
Addr <= "0111010010110";
Trees_din <= "00000100000000000110010000000100";
wait for Clk_period;
Addr <= "0111010010111";
Trees_din <= "00000000000101010011101010000001";
wait for Clk_period;
Addr <= "0111010011000";
Trees_din <= "00000000001001100011101010000001";
wait for Clk_period;
Addr <= "0111010011001";
Trees_din <= "00000011000000000110000100001000";
wait for Clk_period;
Addr <= "0111010011010";
Trees_din <= "00000101000000000011010000000100";
wait for Clk_period;
Addr <= "0111010011011";
Trees_din <= "00000000010000000011101010000001";
wait for Clk_period;
Addr <= "0111010011100";
Trees_din <= "00000000001101100011101010000001";
wait for Clk_period;
Addr <= "0111010011101";
Trees_din <= "00000010000000000000100000000100";
wait for Clk_period;
Addr <= "0111010011110";
Trees_din <= "00000000001110110011101010000001";
wait for Clk_period;
Addr <= "0111010011111";
Trees_din <= "00000000011000010011101010000001";
wait for Clk_period;



----------tree 29-------------------

Addr <= "0111010100000";
Trees_din <= "00000111000000000100111010000000";
wait for Clk_period;
Addr <= "0111010100001";
Trees_din <= "00000010000000000101111001000000";
wait for Clk_period;
Addr <= "0111010100010";
Trees_din <= "00000011000000000100000100100000";
wait for Clk_period;
Addr <= "0111010100011";
Trees_din <= "00000001000000000001001100010000";
wait for Clk_period;
Addr <= "0111010100100";
Trees_din <= "00000000000000000000010100001000";
wait for Clk_period;
Addr <= "0111010100101";
Trees_din <= "00000101000000000000100100000100";
wait for Clk_period;
Addr <= "0111010100110";
Trees_din <= "00000000000111000011110001111111";
wait for Clk_period;
Addr <= "0111010100111";
Trees_din <= "00000000011001000011110001111111";
wait for Clk_period;
Addr <= "0111010101000";
Trees_din <= "00000010000000000001010100000100";
wait for Clk_period;
Addr <= "0111010101001";
Trees_din <= "00000000010011100011110001111111";
wait for Clk_period;
Addr <= "0111010101010";
Trees_din <= "00000000000110110011110001111111";
wait for Clk_period;
Addr <= "0111010101011";
Trees_din <= "00000000000000000110001000001000";
wait for Clk_period;
Addr <= "0111010101100";
Trees_din <= "00000000000000000001110100000100";
wait for Clk_period;
Addr <= "0111010101101";
Trees_din <= "00000000011000110011110001111111";
wait for Clk_period;
Addr <= "0111010101110";
Trees_din <= "00000000010100000011110001111111";
wait for Clk_period;
Addr <= "0111010101111";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "0111010110000";
Trees_din <= "00000000000100100011110001111111";
wait for Clk_period;
Addr <= "0111010110001";
Trees_din <= "00000000011000110011110001111111";
wait for Clk_period;
Addr <= "0111010110010";
Trees_din <= "00000101000000000010100000010000";
wait for Clk_period;
Addr <= "0111010110011";
Trees_din <= "00000101000000000101100100001000";
wait for Clk_period;
Addr <= "0111010110100";
Trees_din <= "00000111000000000110000100000100";
wait for Clk_period;
Addr <= "0111010110101";
Trees_din <= "00000000000011000011110001111111";
wait for Clk_period;
Addr <= "0111010110110";
Trees_din <= "00000000000101000011110001111111";
wait for Clk_period;
Addr <= "0111010110111";
Trees_din <= "00000011000000000001110100000100";
wait for Clk_period;
Addr <= "0111010111000";
Trees_din <= "00000000001001000011110001111111";
wait for Clk_period;
Addr <= "0111010111001";
Trees_din <= "00000000010000010011110001111111";
wait for Clk_period;
Addr <= "0111010111010";
Trees_din <= "00000110000000000000000000001000";
wait for Clk_period;
Addr <= "0111010111011";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "0111010111100";
Trees_din <= "00000000010000110011110001111111";
wait for Clk_period;
Addr <= "0111010111101";
Trees_din <= "00000000001010000011110001111111";
wait for Clk_period;
Addr <= "0111010111110";
Trees_din <= "00000011000000000010001100000100";
wait for Clk_period;
Addr <= "0111010111111";
Trees_din <= "00000000001100000011110001111111";
wait for Clk_period;
Addr <= "0111011000000";
Trees_din <= "00000000010010100011110001111111";
wait for Clk_period;
Addr <= "0111011000001";
Trees_din <= "00000010000000000010011100100000";
wait for Clk_period;
Addr <= "0111011000010";
Trees_din <= "00000111000000000010000100010000";
wait for Clk_period;
Addr <= "0111011000011";
Trees_din <= "00000001000000000011110000001000";
wait for Clk_period;
Addr <= "0111011000100";
Trees_din <= "00000000000000000010101100000100";
wait for Clk_period;
Addr <= "0111011000101";
Trees_din <= "00000000000011010011110001111111";
wait for Clk_period;
Addr <= "0111011000110";
Trees_din <= "00000000010001010011110001111111";
wait for Clk_period;
Addr <= "0111011000111";
Trees_din <= "00000111000000000010101000000100";
wait for Clk_period;
Addr <= "0111011001000";
Trees_din <= "00000000010100000011110001111111";
wait for Clk_period;
Addr <= "0111011001001";
Trees_din <= "00000000001100010011110001111111";
wait for Clk_period;
Addr <= "0111011001010";
Trees_din <= "00000101000000000000000000001000";
wait for Clk_period;
Addr <= "0111011001011";
Trees_din <= "00000010000000000011001100000100";
wait for Clk_period;
Addr <= "0111011001100";
Trees_din <= "00000000001010000011110001111111";
wait for Clk_period;
Addr <= "0111011001101";
Trees_din <= "00000000010101110011110001111111";
wait for Clk_period;
Addr <= "0111011001110";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "0111011001111";
Trees_din <= "00000000000011100011110001111111";
wait for Clk_period;
Addr <= "0111011010000";
Trees_din <= "00000000000000100011110001111111";
wait for Clk_period;
Addr <= "0111011010001";
Trees_din <= "00000110000000000110001100010000";
wait for Clk_period;
Addr <= "0111011010010";
Trees_din <= "00000101000000000011100100001000";
wait for Clk_period;
Addr <= "0111011010011";
Trees_din <= "00000111000000000000101000000100";
wait for Clk_period;
Addr <= "0111011010100";
Trees_din <= "00000000001010000011110001111111";
wait for Clk_period;
Addr <= "0111011010101";
Trees_din <= "00000000000101110011110001111111";
wait for Clk_period;
Addr <= "0111011010110";
Trees_din <= "00000111000000000101000100000100";
wait for Clk_period;
Addr <= "0111011010111";
Trees_din <= "00000000000110110011110001111111";
wait for Clk_period;
Addr <= "0111011011000";
Trees_din <= "00000000000001100011110001111111";
wait for Clk_period;
Addr <= "0111011011001";
Trees_din <= "00000010000000000000000100001000";
wait for Clk_period;
Addr <= "0111011011010";
Trees_din <= "00000111000000000010110100000100";
wait for Clk_period;
Addr <= "0111011011011";
Trees_din <= "00000000001110010011110001111111";
wait for Clk_period;
Addr <= "0111011011100";
Trees_din <= "00000000001010000011110001111111";
wait for Clk_period;
Addr <= "0111011011101";
Trees_din <= "00000101000000000100111100000100";
wait for Clk_period;
Addr <= "0111011011110";
Trees_din <= "00000000001000110011110001111111";
wait for Clk_period;
Addr <= "0111011011111";
Trees_din <= "00000000010111110011110001111111";
wait for Clk_period;
Addr <= "0111011100000";
Trees_din <= "00000101000000000101010101000000";
wait for Clk_period;
Addr <= "0111011100001";
Trees_din <= "00000100000000000010111100100000";
wait for Clk_period;
Addr <= "0111011100010";
Trees_din <= "00000010000000000010011100010000";
wait for Clk_period;
Addr <= "0111011100011";
Trees_din <= "00000110000000000000001100001000";
wait for Clk_period;
Addr <= "0111011100100";
Trees_din <= "00000100000000000101000100000100";
wait for Clk_period;
Addr <= "0111011100101";
Trees_din <= "00000000000101000011110001111111";
wait for Clk_period;
Addr <= "0111011100110";
Trees_din <= "00000000001101000011110001111111";
wait for Clk_period;
Addr <= "0111011100111";
Trees_din <= "00000000000000000001100100000100";
wait for Clk_period;
Addr <= "0111011101000";
Trees_din <= "00000000010000100011110001111111";
wait for Clk_period;
Addr <= "0111011101001";
Trees_din <= "00000000000100010011110001111111";
wait for Clk_period;
Addr <= "0111011101010";
Trees_din <= "00000011000000000000010100001000";
wait for Clk_period;
Addr <= "0111011101011";
Trees_din <= "00000100000000000100001000000100";
wait for Clk_period;
Addr <= "0111011101100";
Trees_din <= "00000000011000000011110001111111";
wait for Clk_period;
Addr <= "0111011101101";
Trees_din <= "00000000010010100011110001111111";
wait for Clk_period;
Addr <= "0111011101110";
Trees_din <= "00000011000000000011111100000100";
wait for Clk_period;
Addr <= "0111011101111";
Trees_din <= "00000000001011010011110001111111";
wait for Clk_period;
Addr <= "0111011110000";
Trees_din <= "00000000010011000011110001111111";
wait for Clk_period;
Addr <= "0111011110001";
Trees_din <= "00000100000000000010100100010000";
wait for Clk_period;
Addr <= "0111011110010";
Trees_din <= "00000001000000000011100100001000";
wait for Clk_period;
Addr <= "0111011110011";
Trees_din <= "00000110000000000010011000000100";
wait for Clk_period;
Addr <= "0111011110100";
Trees_din <= "00000000011000000011110001111111";
wait for Clk_period;
Addr <= "0111011110101";
Trees_din <= "00000000010000100011110001111111";
wait for Clk_period;
Addr <= "0111011110110";
Trees_din <= "00000011000000000011110100000100";
wait for Clk_period;
Addr <= "0111011110111";
Trees_din <= "00000000000100100011110001111111";
wait for Clk_period;
Addr <= "0111011111000";
Trees_din <= "00000000001110110011110001111111";
wait for Clk_period;
Addr <= "0111011111001";
Trees_din <= "00000001000000000011100000001000";
wait for Clk_period;
Addr <= "0111011111010";
Trees_din <= "00000110000000000001101000000100";
wait for Clk_period;
Addr <= "0111011111011";
Trees_din <= "00000000000111100011110001111111";
wait for Clk_period;
Addr <= "0111011111100";
Trees_din <= "00000000010111000011110001111111";
wait for Clk_period;
Addr <= "0111011111101";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "0111011111110";
Trees_din <= "00000000000001100011110001111111";
wait for Clk_period;
Addr <= "0111011111111";
Trees_din <= "00000000000110110011110001111111";
wait for Clk_period;
Addr <= "0111100000000";
Trees_din <= "00000110000000000000100100100000";
wait for Clk_period;
Addr <= "0111100000001";
Trees_din <= "00000101000000000101000000010000";
wait for Clk_period;
Addr <= "0111100000010";
Trees_din <= "00000000000000000100110000001000";
wait for Clk_period;
Addr <= "0111100000011";
Trees_din <= "00000101000000000100100000000100";
wait for Clk_period;
Addr <= "0111100000100";
Trees_din <= "00000000001010100011110001111111";
wait for Clk_period;
Addr <= "0111100000101";
Trees_din <= "00000000000011100011110001111111";
wait for Clk_period;
Addr <= "0111100000110";
Trees_din <= "00000000000000000000110000000100";
wait for Clk_period;
Addr <= "0111100000111";
Trees_din <= "00000000010011010011110001111111";
wait for Clk_period;
Addr <= "0111100001000";
Trees_din <= "00000000000110000011110001111111";
wait for Clk_period;
Addr <= "0111100001001";
Trees_din <= "00000110000000000100110100001000";
wait for Clk_period;
Addr <= "0111100001010";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "0111100001011";
Trees_din <= "00000000001001100011110001111111";
wait for Clk_period;
Addr <= "0111100001100";
Trees_din <= "00000000001101100011110001111111";
wait for Clk_period;
Addr <= "0111100001101";
Trees_din <= "00000101000000000010100100000100";
wait for Clk_period;
Addr <= "0111100001110";
Trees_din <= "00000000010001100011110001111111";
wait for Clk_period;
Addr <= "0111100001111";
Trees_din <= "00000000001001100011110001111111";
wait for Clk_period;
Addr <= "0111100010000";
Trees_din <= "00000100000000000101000000010000";
wait for Clk_period;
Addr <= "0111100010001";
Trees_din <= "00000101000000000011010000001000";
wait for Clk_period;
Addr <= "0111100010010";
Trees_din <= "00000001000000000011110000000100";
wait for Clk_period;
Addr <= "0111100010011";
Trees_din <= "00000000011000000011110001111111";
wait for Clk_period;
Addr <= "0111100010100";
Trees_din <= "00000000000100100011110001111111";
wait for Clk_period;
Addr <= "0111100010101";
Trees_din <= "00000010000000000000000100000100";
wait for Clk_period;
Addr <= "0111100010110";
Trees_din <= "00000000000011000011110001111111";
wait for Clk_period;
Addr <= "0111100010111";
Trees_din <= "00000000010110110011110001111111";
wait for Clk_period;
Addr <= "0111100011000";
Trees_din <= "00000100000000000100011100001000";
wait for Clk_period;
Addr <= "0111100011001";
Trees_din <= "00000001000000000011000100000100";
wait for Clk_period;
Addr <= "0111100011010";
Trees_din <= "00000000000000010011110001111111";
wait for Clk_period;
Addr <= "0111100011011";
Trees_din <= "00000000000001010011110001111111";
wait for Clk_period;
Addr <= "0111100011100";
Trees_din <= "00000011000000000011011000000100";
wait for Clk_period;
Addr <= "0111100011101";
Trees_din <= "00000000010011010011110001111111";
wait for Clk_period;
Addr <= "0111100011110";
Trees_din <= "00000000000101010011110001111111";
wait for Clk_period;



----------tree 30-------------------

Addr <= "0111100011111";
Trees_din <= "00000110000000000010111010000000";
wait for Clk_period;
Addr <= "0111100100000";
Trees_din <= "00000000000000000000100101000000";
wait for Clk_period;
Addr <= "0111100100001";
Trees_din <= "00000101000000000100010000100000";
wait for Clk_period;
Addr <= "0111100100010";
Trees_din <= "00000010000000000010010000010000";
wait for Clk_period;
Addr <= "0111100100011";
Trees_din <= "00000101000000000001000000001000";
wait for Clk_period;
Addr <= "0111100100100";
Trees_din <= "00000100000000000010010100000100";
wait for Clk_period;
Addr <= "0111100100101";
Trees_din <= "00000000010101110011111001111001";
wait for Clk_period;
Addr <= "0111100100110";
Trees_din <= "00000000010011110011111001111001";
wait for Clk_period;
Addr <= "0111100100111";
Trees_din <= "00000110000000000101000000000100";
wait for Clk_period;
Addr <= "0111100101000";
Trees_din <= "00000000000111000011111001111001";
wait for Clk_period;
Addr <= "0111100101001";
Trees_din <= "00000000001010100011111001111001";
wait for Clk_period;
Addr <= "0111100101010";
Trees_din <= "00000111000000000000011100001000";
wait for Clk_period;
Addr <= "0111100101011";
Trees_din <= "00000001000000000101000000000100";
wait for Clk_period;
Addr <= "0111100101100";
Trees_din <= "00000000001010100011111001111001";
wait for Clk_period;
Addr <= "0111100101101";
Trees_din <= "00000000000001000011111001111001";
wait for Clk_period;
Addr <= "0111100101110";
Trees_din <= "00000110000000000100100100000100";
wait for Clk_period;
Addr <= "0111100101111";
Trees_din <= "00000000010001110011111001111001";
wait for Clk_period;
Addr <= "0111100110000";
Trees_din <= "00000000001001000011111001111001";
wait for Clk_period;
Addr <= "0111100110001";
Trees_din <= "00000111000000000110001000010000";
wait for Clk_period;
Addr <= "0111100110010";
Trees_din <= "00000101000000000110001000001000";
wait for Clk_period;
Addr <= "0111100110011";
Trees_din <= "00000001000000000001000000000100";
wait for Clk_period;
Addr <= "0111100110100";
Trees_din <= "00000000010100110011111001111001";
wait for Clk_period;
Addr <= "0111100110101";
Trees_din <= "00000000001010100011111001111001";
wait for Clk_period;
Addr <= "0111100110110";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "0111100110111";
Trees_din <= "00000000000100000011111001111001";
wait for Clk_period;
Addr <= "0111100111000";
Trees_din <= "00000000001101110011111001111001";
wait for Clk_period;
Addr <= "0111100111001";
Trees_din <= "00000000000000000100111000001000";
wait for Clk_period;
Addr <= "0111100111010";
Trees_din <= "00000000000000000010011100000100";
wait for Clk_period;
Addr <= "0111100111011";
Trees_din <= "00000000011001000011111001111001";
wait for Clk_period;
Addr <= "0111100111100";
Trees_din <= "00000000001001110011111001111001";
wait for Clk_period;
Addr <= "0111100111101";
Trees_din <= "00000000000000000010101000000100";
wait for Clk_period;
Addr <= "0111100111110";
Trees_din <= "00000000000000100011111001111001";
wait for Clk_period;
Addr <= "0111100111111";
Trees_din <= "00000000001101000011111001111001";
wait for Clk_period;
Addr <= "0111101000000";
Trees_din <= "00000001000000000100101100100000";
wait for Clk_period;
Addr <= "0111101000001";
Trees_din <= "00000010000000000000101000010000";
wait for Clk_period;
Addr <= "0111101000010";
Trees_din <= "00000110000000000101100000001000";
wait for Clk_period;
Addr <= "0111101000011";
Trees_din <= "00000101000000000000110100000100";
wait for Clk_period;
Addr <= "0111101000100";
Trees_din <= "00000000000000010011111001111001";
wait for Clk_period;
Addr <= "0111101000101";
Trees_din <= "00000000010000100011111001111001";
wait for Clk_period;
Addr <= "0111101000110";
Trees_din <= "00000101000000000011001100000100";
wait for Clk_period;
Addr <= "0111101000111";
Trees_din <= "00000000000110010011111001111001";
wait for Clk_period;
Addr <= "0111101001000";
Trees_din <= "00000000001010000011111001111001";
wait for Clk_period;
Addr <= "0111101001001";
Trees_din <= "00000011000000000100001000001000";
wait for Clk_period;
Addr <= "0111101001010";
Trees_din <= "00000101000000000100001000000100";
wait for Clk_period;
Addr <= "0111101001011";
Trees_din <= "00000000010010110011111001111001";
wait for Clk_period;
Addr <= "0111101001100";
Trees_din <= "00000000010101010011111001111001";
wait for Clk_period;
Addr <= "0111101001101";
Trees_din <= "00000011000000000100100100000100";
wait for Clk_period;
Addr <= "0111101001110";
Trees_din <= "00000000000110000011111001111001";
wait for Clk_period;
Addr <= "0111101001111";
Trees_din <= "00000000000100010011111001111001";
wait for Clk_period;
Addr <= "0111101010000";
Trees_din <= "00000111000000000011100100010000";
wait for Clk_period;
Addr <= "0111101010001";
Trees_din <= "00000011000000000011100000001000";
wait for Clk_period;
Addr <= "0111101010010";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "0111101010011";
Trees_din <= "00000000001100100011111001111001";
wait for Clk_period;
Addr <= "0111101010100";
Trees_din <= "00000000001100000011111001111001";
wait for Clk_period;
Addr <= "0111101010101";
Trees_din <= "00000011000000000001111000000100";
wait for Clk_period;
Addr <= "0111101010110";
Trees_din <= "00000000001010100011111001111001";
wait for Clk_period;
Addr <= "0111101010111";
Trees_din <= "00000000010110110011111001111001";
wait for Clk_period;
Addr <= "0111101011000";
Trees_din <= "00000100000000000100110000001000";
wait for Clk_period;
Addr <= "0111101011001";
Trees_din <= "00000101000000000100001100000100";
wait for Clk_period;
Addr <= "0111101011010";
Trees_din <= "00000000000001000011111001111001";
wait for Clk_period;
Addr <= "0111101011011";
Trees_din <= "00000000010011010011111001111001";
wait for Clk_period;
Addr <= "0111101011100";
Trees_din <= "00000000000000000010000000000100";
wait for Clk_period;
Addr <= "0111101011101";
Trees_din <= "00000000001011010011111001111001";
wait for Clk_period;
Addr <= "0111101011110";
Trees_din <= "00000000001111000011111001111001";
wait for Clk_period;
Addr <= "0111101011111";
Trees_din <= "00000110000000000011000101000000";
wait for Clk_period;
Addr <= "0111101100000";
Trees_din <= "00000111000000000101110100100000";
wait for Clk_period;
Addr <= "0111101100001";
Trees_din <= "00000100000000000011010000010000";
wait for Clk_period;
Addr <= "0111101100010";
Trees_din <= "00000011000000000101110100001000";
wait for Clk_period;
Addr <= "0111101100011";
Trees_din <= "00000001000000000101001000000100";
wait for Clk_period;
Addr <= "0111101100100";
Trees_din <= "00000000010110110011111001111001";
wait for Clk_period;
Addr <= "0111101100101";
Trees_din <= "00000000000011110011111001111001";
wait for Clk_period;
Addr <= "0111101100110";
Trees_din <= "00000101000000000100000100000100";
wait for Clk_period;
Addr <= "0111101100111";
Trees_din <= "00000000010001010011111001111001";
wait for Clk_period;
Addr <= "0111101101000";
Trees_din <= "00000000001100000011111001111001";
wait for Clk_period;
Addr <= "0111101101001";
Trees_din <= "00000101000000000011100100001000";
wait for Clk_period;
Addr <= "0111101101010";
Trees_din <= "00000111000000000101010100000100";
wait for Clk_period;
Addr <= "0111101101011";
Trees_din <= "00000000000001110011111001111001";
wait for Clk_period;
Addr <= "0111101101100";
Trees_din <= "00000000000100000011111001111001";
wait for Clk_period;
Addr <= "0111101101101";
Trees_din <= "00000100000000000000110100000100";
wait for Clk_period;
Addr <= "0111101101110";
Trees_din <= "00000000000000100011111001111001";
wait for Clk_period;
Addr <= "0111101101111";
Trees_din <= "00000000011000110011111001111001";
wait for Clk_period;
Addr <= "0111101110000";
Trees_din <= "00000001000000000011011100010000";
wait for Clk_period;
Addr <= "0111101110001";
Trees_din <= "00000111000000000000100000001000";
wait for Clk_period;
Addr <= "0111101110010";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "0111101110011";
Trees_din <= "00000000001001100011111001111001";
wait for Clk_period;
Addr <= "0111101110100";
Trees_din <= "00000000001001100011111001111001";
wait for Clk_period;
Addr <= "0111101110101";
Trees_din <= "00000000000000000011110000000100";
wait for Clk_period;
Addr <= "0111101110110";
Trees_din <= "00000000001010110011111001111001";
wait for Clk_period;
Addr <= "0111101110111";
Trees_din <= "00000000001111000011111001111001";
wait for Clk_period;
Addr <= "0111101111000";
Trees_din <= "00000100000000000000101100001000";
wait for Clk_period;
Addr <= "0111101111001";
Trees_din <= "00000111000000000101100100000100";
wait for Clk_period;
Addr <= "0111101111010";
Trees_din <= "00000000000101110011111001111001";
wait for Clk_period;
Addr <= "0111101111011";
Trees_din <= "00000000010100100011111001111001";
wait for Clk_period;
Addr <= "0111101111100";
Trees_din <= "00000111000000000011100100000100";
wait for Clk_period;
Addr <= "0111101111101";
Trees_din <= "00000000000100000011111001111001";
wait for Clk_period;
Addr <= "0111101111110";
Trees_din <= "00000000010110000011111001111001";
wait for Clk_period;
Addr <= "0111101111111";
Trees_din <= "00000111000000000011000100100000";
wait for Clk_period;
Addr <= "0111110000000";
Trees_din <= "00000110000000000110001100010000";
wait for Clk_period;
Addr <= "0111110000001";
Trees_din <= "00000110000000000001111000001000";
wait for Clk_period;
Addr <= "0111110000010";
Trees_din <= "00000111000000000000000000000100";
wait for Clk_period;
Addr <= "0111110000011";
Trees_din <= "00000000010011110011111001111001";
wait for Clk_period;
Addr <= "0111110000100";
Trees_din <= "00000000001001100011111001111001";
wait for Clk_period;
Addr <= "0111110000101";
Trees_din <= "00000001000000000100100000000100";
wait for Clk_period;
Addr <= "0111110000110";
Trees_din <= "00000000010101110011111001111001";
wait for Clk_period;
Addr <= "0111110000111";
Trees_din <= "00000000000011010011111001111001";
wait for Clk_period;
Addr <= "0111110001000";
Trees_din <= "00000100000000000101111000001000";
wait for Clk_period;
Addr <= "0111110001001";
Trees_din <= "00000001000000000010100100000100";
wait for Clk_period;
Addr <= "0111110001010";
Trees_din <= "00000000001110110011111001111001";
wait for Clk_period;
Addr <= "0111110001011";
Trees_din <= "00000000010101100011111001111001";
wait for Clk_period;
Addr <= "0111110001100";
Trees_din <= "00000010000000000000001000000100";
wait for Clk_period;
Addr <= "0111110001101";
Trees_din <= "00000000010000100011111001111001";
wait for Clk_period;
Addr <= "0111110001110";
Trees_din <= "00000000001000110011111001111001";
wait for Clk_period;
Addr <= "0111110001111";
Trees_din <= "00000001000000000010011100010000";
wait for Clk_period;
Addr <= "0111110010000";
Trees_din <= "00000001000000000101110000001000";
wait for Clk_period;
Addr <= "0111110010001";
Trees_din <= "00000110000000000010010100000100";
wait for Clk_period;
Addr <= "0111110010010";
Trees_din <= "00000000010010010011111001111001";
wait for Clk_period;
Addr <= "0111110010011";
Trees_din <= "00000000010011000011111001111001";
wait for Clk_period;
Addr <= "0111110010100";
Trees_din <= "00000111000000000100110100000100";
wait for Clk_period;
Addr <= "0111110010101";
Trees_din <= "00000000010110110011111001111001";
wait for Clk_period;
Addr <= "0111110010110";
Trees_din <= "00000000001001100011111001111001";
wait for Clk_period;
Addr <= "0111110010111";
Trees_din <= "00000101000000000100010100001000";
wait for Clk_period;
Addr <= "0111110011000";
Trees_din <= "00000110000000000001010000000100";
wait for Clk_period;
Addr <= "0111110011001";
Trees_din <= "00000000001111010011111001111001";
wait for Clk_period;
Addr <= "0111110011010";
Trees_din <= "00000000011000010011111001111001";
wait for Clk_period;
Addr <= "0111110011011";
Trees_din <= "00000011000000000010101100000100";
wait for Clk_period;
Addr <= "0111110011100";
Trees_din <= "00000000010001100011111001111001";
wait for Clk_period;
Addr <= "0111110011101";
Trees_din <= "00000000010110010011111001111001";
wait for Clk_period;



----------tree 31-------------------

Addr <= "0111110011110";
Trees_din <= "00000100000000000101010010000000";
wait for Clk_period;
Addr <= "0111110011111";
Trees_din <= "00000100000000000001010001000000";
wait for Clk_period;
Addr <= "0111110100000";
Trees_din <= "00000011000000000101100100100000";
wait for Clk_period;
Addr <= "0111110100001";
Trees_din <= "00000111000000000011001100010000";
wait for Clk_period;
Addr <= "0111110100010";
Trees_din <= "00000100000000000001010000001000";
wait for Clk_period;
Addr <= "0111110100011";
Trees_din <= "00000100000000000101100000000100";
wait for Clk_period;
Addr <= "0111110100100";
Trees_din <= "00000000000001000100000001110101";
wait for Clk_period;
Addr <= "0111110100101";
Trees_din <= "00000000001101110100000001110101";
wait for Clk_period;
Addr <= "0111110100110";
Trees_din <= "00000111000000000000000100000100";
wait for Clk_period;
Addr <= "0111110100111";
Trees_din <= "00000000000010110100000001110101";
wait for Clk_period;
Addr <= "0111110101000";
Trees_din <= "00000000000001010100000001110101";
wait for Clk_period;
Addr <= "0111110101001";
Trees_din <= "00000101000000000000011000001000";
wait for Clk_period;
Addr <= "0111110101010";
Trees_din <= "00000010000000000001101100000100";
wait for Clk_period;
Addr <= "0111110101011";
Trees_din <= "00000000001100010100000001110101";
wait for Clk_period;
Addr <= "0111110101100";
Trees_din <= "00000000001100000100000001110101";
wait for Clk_period;
Addr <= "0111110101101";
Trees_din <= "00000001000000000001110000000100";
wait for Clk_period;
Addr <= "0111110101110";
Trees_din <= "00000000001000100100000001110101";
wait for Clk_period;
Addr <= "0111110101111";
Trees_din <= "00000000000000100100000001110101";
wait for Clk_period;
Addr <= "0111110110000";
Trees_din <= "00000010000000000101010000010000";
wait for Clk_period;
Addr <= "0111110110001";
Trees_din <= "00000001000000000100010100001000";
wait for Clk_period;
Addr <= "0111110110010";
Trees_din <= "00000110000000000011111100000100";
wait for Clk_period;
Addr <= "0111110110011";
Trees_din <= "00000000001011010100000001110101";
wait for Clk_period;
Addr <= "0111110110100";
Trees_din <= "00000000011000000100000001110101";
wait for Clk_period;
Addr <= "0111110110101";
Trees_din <= "00000110000000000011101100000100";
wait for Clk_period;
Addr <= "0111110110110";
Trees_din <= "00000000011000110100000001110101";
wait for Clk_period;
Addr <= "0111110110111";
Trees_din <= "00000000000010110100000001110101";
wait for Clk_period;
Addr <= "0111110111000";
Trees_din <= "00000100000000000100001100001000";
wait for Clk_period;
Addr <= "0111110111001";
Trees_din <= "00000000000000000100101100000100";
wait for Clk_period;
Addr <= "0111110111010";
Trees_din <= "00000000010011010100000001110101";
wait for Clk_period;
Addr <= "0111110111011";
Trees_din <= "00000000000111100100000001110101";
wait for Clk_period;
Addr <= "0111110111100";
Trees_din <= "00000001000000000100111000000100";
wait for Clk_period;
Addr <= "0111110111101";
Trees_din <= "00000000010010010100000001110101";
wait for Clk_period;
Addr <= "0111110111110";
Trees_din <= "00000000001101110100000001110101";
wait for Clk_period;
Addr <= "0111110111111";
Trees_din <= "00000110000000000001100100100000";
wait for Clk_period;
Addr <= "0111111000000";
Trees_din <= "00000110000000000000000000010000";
wait for Clk_period;
Addr <= "0111111000001";
Trees_din <= "00000110000000000101001000001000";
wait for Clk_period;
Addr <= "0111111000010";
Trees_din <= "00000011000000000000101000000100";
wait for Clk_period;
Addr <= "0111111000011";
Trees_din <= "00000000010110000100000001110101";
wait for Clk_period;
Addr <= "0111111000100";
Trees_din <= "00000000010000010100000001110101";
wait for Clk_period;
Addr <= "0111111000101";
Trees_din <= "00000011000000000011100000000100";
wait for Clk_period;
Addr <= "0111111000110";
Trees_din <= "00000000010010100100000001110101";
wait for Clk_period;
Addr <= "0111111000111";
Trees_din <= "00000000001011100100000001110101";
wait for Clk_period;
Addr <= "0111111001000";
Trees_din <= "00000101000000000100010100001000";
wait for Clk_period;
Addr <= "0111111001001";
Trees_din <= "00000001000000000000010100000100";
wait for Clk_period;
Addr <= "0111111001010";
Trees_din <= "00000000001001100100000001110101";
wait for Clk_period;
Addr <= "0111111001011";
Trees_din <= "00000000000010010100000001110101";
wait for Clk_period;
Addr <= "0111111001100";
Trees_din <= "00000101000000000101110000000100";
wait for Clk_period;
Addr <= "0111111001101";
Trees_din <= "00000000010011010100000001110101";
wait for Clk_period;
Addr <= "0111111001110";
Trees_din <= "00000000001011110100000001110101";
wait for Clk_period;
Addr <= "0111111001111";
Trees_din <= "00000110000000000010000100010000";
wait for Clk_period;
Addr <= "0111111010000";
Trees_din <= "00000001000000000011001100001000";
wait for Clk_period;
Addr <= "0111111010001";
Trees_din <= "00000010000000000100100000000100";
wait for Clk_period;
Addr <= "0111111010010";
Trees_din <= "00000000001001100100000001110101";
wait for Clk_period;
Addr <= "0111111010011";
Trees_din <= "00000000001011010100000001110101";
wait for Clk_period;
Addr <= "0111111010100";
Trees_din <= "00000010000000000000010100000100";
wait for Clk_period;
Addr <= "0111111010101";
Trees_din <= "00000000000100110100000001110101";
wait for Clk_period;
Addr <= "0111111010110";
Trees_din <= "00000000000101010100000001110101";
wait for Clk_period;
Addr <= "0111111010111";
Trees_din <= "00000101000000000000110000001000";
wait for Clk_period;
Addr <= "0111111011000";
Trees_din <= "00000001000000000010011100000100";
wait for Clk_period;
Addr <= "0111111011001";
Trees_din <= "00000000000010010100000001110101";
wait for Clk_period;
Addr <= "0111111011010";
Trees_din <= "00000000000101000100000001110101";
wait for Clk_period;
Addr <= "0111111011011";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "0111111011100";
Trees_din <= "00000000001010100100000001110101";
wait for Clk_period;
Addr <= "0111111011101";
Trees_din <= "00000000001100000100000001110101";
wait for Clk_period;
Addr <= "0111111011110";
Trees_din <= "00000101000000000001001001000000";
wait for Clk_period;
Addr <= "0111111011111";
Trees_din <= "00000001000000000001010000100000";
wait for Clk_period;
Addr <= "0111111100000";
Trees_din <= "00000100000000000001000000010000";
wait for Clk_period;
Addr <= "0111111100001";
Trees_din <= "00000100000000000001010100001000";
wait for Clk_period;
Addr <= "0111111100010";
Trees_din <= "00000000000000000101001000000100";
wait for Clk_period;
Addr <= "0111111100011";
Trees_din <= "00000000010110000100000001110101";
wait for Clk_period;
Addr <= "0111111100100";
Trees_din <= "00000000000000100100000001110101";
wait for Clk_period;
Addr <= "0111111100101";
Trees_din <= "00000001000000000011110100000100";
wait for Clk_period;
Addr <= "0111111100110";
Trees_din <= "00000000000001100100000001110101";
wait for Clk_period;
Addr <= "0111111100111";
Trees_din <= "00000000010001000100000001110101";
wait for Clk_period;
Addr <= "0111111101000";
Trees_din <= "00000111000000000000101000001000";
wait for Clk_period;
Addr <= "0111111101001";
Trees_din <= "00000111000000000101101000000100";
wait for Clk_period;
Addr <= "0111111101010";
Trees_din <= "00000000011001000100000001110101";
wait for Clk_period;
Addr <= "0111111101011";
Trees_din <= "00000000010111010100000001110101";
wait for Clk_period;
Addr <= "0111111101100";
Trees_din <= "00000011000000000101000000000100";
wait for Clk_period;
Addr <= "0111111101101";
Trees_din <= "00000000010010010100000001110101";
wait for Clk_period;
Addr <= "0111111101110";
Trees_din <= "00000000001001010100000001110101";
wait for Clk_period;
Addr <= "0111111101111";
Trees_din <= "00000010000000000010010000010000";
wait for Clk_period;
Addr <= "0111111110000";
Trees_din <= "00000100000000000000000000001000";
wait for Clk_period;
Addr <= "0111111110001";
Trees_din <= "00000101000000000010001000000100";
wait for Clk_period;
Addr <= "0111111110010";
Trees_din <= "00000000010011110100000001110101";
wait for Clk_period;
Addr <= "0111111110011";
Trees_din <= "00000000001100110100000001110101";
wait for Clk_period;
Addr <= "0111111110100";
Trees_din <= "00000011000000000010101100000100";
wait for Clk_period;
Addr <= "0111111110101";
Trees_din <= "00000000011000110100000001110101";
wait for Clk_period;
Addr <= "0111111110110";
Trees_din <= "00000000010011100100000001110101";
wait for Clk_period;
Addr <= "0111111110111";
Trees_din <= "00000011000000000100010100001000";
wait for Clk_period;
Addr <= "0111111111000";
Trees_din <= "00000110000000000001111100000100";
wait for Clk_period;
Addr <= "0111111111001";
Trees_din <= "00000000010101000100000001110101";
wait for Clk_period;
Addr <= "0111111111010";
Trees_din <= "00000000000111010100000001110101";
wait for Clk_period;
Addr <= "0111111111011";
Trees_din <= "00000010000000000011110100000100";
wait for Clk_period;
Addr <= "0111111111100";
Trees_din <= "00000000010100010100000001110101";
wait for Clk_period;
Addr <= "0111111111101";
Trees_din <= "00000000010100010100000001110101";
wait for Clk_period;
Addr <= "0111111111110";
Trees_din <= "00000011000000000011110100100000";
wait for Clk_period;
Addr <= "0111111111111";
Trees_din <= "00000001000000000001111000010000";
wait for Clk_period;
Addr <= "1000000000000";
Trees_din <= "00000111000000000101110100001000";
wait for Clk_period;
Addr <= "1000000000001";
Trees_din <= "00000101000000000000010100000100";
wait for Clk_period;
Addr <= "1000000000010";
Trees_din <= "00000000000110000100000001110101";
wait for Clk_period;
Addr <= "1000000000011";
Trees_din <= "00000000000001010100000001110101";
wait for Clk_period;
Addr <= "1000000000100";
Trees_din <= "00000101000000000011011000000100";
wait for Clk_period;
Addr <= "1000000000101";
Trees_din <= "00000000001011110100000001110101";
wait for Clk_period;
Addr <= "1000000000110";
Trees_din <= "00000000010101000100000001110101";
wait for Clk_period;
Addr <= "1000000000111";
Trees_din <= "00000011000000000001101100001000";
wait for Clk_period;
Addr <= "1000000001000";
Trees_din <= "00000100000000000000001100000100";
wait for Clk_period;
Addr <= "1000000001001";
Trees_din <= "00000000000011000100000001110101";
wait for Clk_period;
Addr <= "1000000001010";
Trees_din <= "00000000010010000100000001110101";
wait for Clk_period;
Addr <= "1000000001011";
Trees_din <= "00000001000000000110010000000100";
wait for Clk_period;
Addr <= "1000000001100";
Trees_din <= "00000000001010100100000001110101";
wait for Clk_period;
Addr <= "1000000001101";
Trees_din <= "00000000000100010100000001110101";
wait for Clk_period;
Addr <= "1000000001110";
Trees_din <= "00000001000000000000100000010000";
wait for Clk_period;
Addr <= "1000000001111";
Trees_din <= "00000001000000000011110100001000";
wait for Clk_period;
Addr <= "1000000010000";
Trees_din <= "00000101000000000010100100000100";
wait for Clk_period;
Addr <= "1000000010001";
Trees_din <= "00000000010110110100000001110101";
wait for Clk_period;
Addr <= "1000000010010";
Trees_din <= "00000000000111000100000001110101";
wait for Clk_period;
Addr <= "1000000010011";
Trees_din <= "00000100000000000010001000000100";
wait for Clk_period;
Addr <= "1000000010100";
Trees_din <= "00000000000101100100000001110101";
wait for Clk_period;
Addr <= "1000000010101";
Trees_din <= "00000000000010100100000001110101";
wait for Clk_period;
Addr <= "1000000010110";
Trees_din <= "00000010000000000101101000001000";
wait for Clk_period;
Addr <= "1000000010111";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "1000000011000";
Trees_din <= "00000000000000000100000001110101";
wait for Clk_period;
Addr <= "1000000011001";
Trees_din <= "00000000011000100100000001110101";
wait for Clk_period;
Addr <= "1000000011010";
Trees_din <= "00000111000000000101011000000100";
wait for Clk_period;
Addr <= "1000000011011";
Trees_din <= "00000000001010100100000001110101";
wait for Clk_period;
Addr <= "1000000011100";
Trees_din <= "00000000001110100100000001110101";
wait for Clk_period;



----------tree 32-------------------

Addr <= "1000000011101";
Trees_din <= "00000001000000000101011010000000";
wait for Clk_period;
Addr <= "1000000011110";
Trees_din <= "00000111000000000011111001000000";
wait for Clk_period;
Addr <= "1000000011111";
Trees_din <= "00000101000000000010111100100000";
wait for Clk_period;
Addr <= "1000000100000";
Trees_din <= "00000000000000000010110100010000";
wait for Clk_period;
Addr <= "1000000100001";
Trees_din <= "00000000000000000010100000001000";
wait for Clk_period;
Addr <= "1000000100010";
Trees_din <= "00000000000000000100010100000100";
wait for Clk_period;
Addr <= "1000000100011";
Trees_din <= "00000000001001010100001001110001";
wait for Clk_period;
Addr <= "1000000100100";
Trees_din <= "00000000000001100100001001110001";
wait for Clk_period;
Addr <= "1000000100101";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "1000000100110";
Trees_din <= "00000000001011000100001001110001";
wait for Clk_period;
Addr <= "1000000100111";
Trees_din <= "00000000011000110100001001110001";
wait for Clk_period;
Addr <= "1000000101000";
Trees_din <= "00000010000000000001011100001000";
wait for Clk_period;
Addr <= "1000000101001";
Trees_din <= "00000000000000000011000000000100";
wait for Clk_period;
Addr <= "1000000101010";
Trees_din <= "00000000001011010100001001110001";
wait for Clk_period;
Addr <= "1000000101011";
Trees_din <= "00000000000011100100001001110001";
wait for Clk_period;
Addr <= "1000000101100";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "1000000101101";
Trees_din <= "00000000000010100100001001110001";
wait for Clk_period;
Addr <= "1000000101110";
Trees_din <= "00000000001101010100001001110001";
wait for Clk_period;
Addr <= "1000000101111";
Trees_din <= "00000011000000000101100100010000";
wait for Clk_period;
Addr <= "1000000110000";
Trees_din <= "00000010000000000011101100001000";
wait for Clk_period;
Addr <= "1000000110001";
Trees_din <= "00000011000000000011110000000100";
wait for Clk_period;
Addr <= "1000000110010";
Trees_din <= "00000000001111000100001001110001";
wait for Clk_period;
Addr <= "1000000110011";
Trees_din <= "00000000010001100100001001110001";
wait for Clk_period;
Addr <= "1000000110100";
Trees_din <= "00000011000000000010110000000100";
wait for Clk_period;
Addr <= "1000000110101";
Trees_din <= "00000000001100100100001001110001";
wait for Clk_period;
Addr <= "1000000110110";
Trees_din <= "00000000001101000100001001110001";
wait for Clk_period;
Addr <= "1000000110111";
Trees_din <= "00000001000000000000111000001000";
wait for Clk_period;
Addr <= "1000000111000";
Trees_din <= "00000111000000000000001100000100";
wait for Clk_period;
Addr <= "1000000111001";
Trees_din <= "00000000000011110100001001110001";
wait for Clk_period;
Addr <= "1000000111010";
Trees_din <= "00000000000110010100001001110001";
wait for Clk_period;
Addr <= "1000000111011";
Trees_din <= "00000100000000000101110100000100";
wait for Clk_period;
Addr <= "1000000111100";
Trees_din <= "00000000000010110100001001110001";
wait for Clk_period;
Addr <= "1000000111101";
Trees_din <= "00000000010100010100001001110001";
wait for Clk_period;
Addr <= "1000000111110";
Trees_din <= "00000010000000000001010000100000";
wait for Clk_period;
Addr <= "1000000111111";
Trees_din <= "00000110000000000101001000010000";
wait for Clk_period;
Addr <= "1000001000000";
Trees_din <= "00000011000000000100001000001000";
wait for Clk_period;
Addr <= "1000001000001";
Trees_din <= "00000111000000000011111000000100";
wait for Clk_period;
Addr <= "1000001000010";
Trees_din <= "00000000010000110100001001110001";
wait for Clk_period;
Addr <= "1000001000011";
Trees_din <= "00000000001000000100001001110001";
wait for Clk_period;
Addr <= "1000001000100";
Trees_din <= "00000001000000000001000000000100";
wait for Clk_period;
Addr <= "1000001000101";
Trees_din <= "00000000010010100100001001110001";
wait for Clk_period;
Addr <= "1000001000110";
Trees_din <= "00000000001001100100001001110001";
wait for Clk_period;
Addr <= "1000001000111";
Trees_din <= "00000000000000000000110100001000";
wait for Clk_period;
Addr <= "1000001001000";
Trees_din <= "00000001000000000000100100000100";
wait for Clk_period;
Addr <= "1000001001001";
Trees_din <= "00000000010100010100001001110001";
wait for Clk_period;
Addr <= "1000001001010";
Trees_din <= "00000000001111100100001001110001";
wait for Clk_period;
Addr <= "1000001001011";
Trees_din <= "00000000000000000000011000000100";
wait for Clk_period;
Addr <= "1000001001100";
Trees_din <= "00000000001000000100001001110001";
wait for Clk_period;
Addr <= "1000001001101";
Trees_din <= "00000000010010100100001001110001";
wait for Clk_period;
Addr <= "1000001001110";
Trees_din <= "00000011000000000010110000010000";
wait for Clk_period;
Addr <= "1000001001111";
Trees_din <= "00000111000000000100111000001000";
wait for Clk_period;
Addr <= "1000001010000";
Trees_din <= "00000101000000000011011100000100";
wait for Clk_period;
Addr <= "1000001010001";
Trees_din <= "00000000000101110100001001110001";
wait for Clk_period;
Addr <= "1000001010010";
Trees_din <= "00000000011000010100001001110001";
wait for Clk_period;
Addr <= "1000001010011";
Trees_din <= "00000000000000000011011000000100";
wait for Clk_period;
Addr <= "1000001010100";
Trees_din <= "00000000010011000100001001110001";
wait for Clk_period;
Addr <= "1000001010101";
Trees_din <= "00000000010111110100001001110001";
wait for Clk_period;
Addr <= "1000001010110";
Trees_din <= "00000001000000000100011100001000";
wait for Clk_period;
Addr <= "1000001010111";
Trees_din <= "00000001000000000100111100000100";
wait for Clk_period;
Addr <= "1000001011000";
Trees_din <= "00000000001110010100001001110001";
wait for Clk_period;
Addr <= "1000001011001";
Trees_din <= "00000000001101110100001001110001";
wait for Clk_period;
Addr <= "1000001011010";
Trees_din <= "00000111000000000010010000000100";
wait for Clk_period;
Addr <= "1000001011011";
Trees_din <= "00000000010100110100001001110001";
wait for Clk_period;
Addr <= "1000001011100";
Trees_din <= "00000000010100110100001001110001";
wait for Clk_period;
Addr <= "1000001011101";
Trees_din <= "00000011000000000101111001000000";
wait for Clk_period;
Addr <= "1000001011110";
Trees_din <= "00000100000000000100110000100000";
wait for Clk_period;
Addr <= "1000001011111";
Trees_din <= "00000100000000000001110000010000";
wait for Clk_period;
Addr <= "1000001100000";
Trees_din <= "00000100000000000001110100001000";
wait for Clk_period;
Addr <= "1000001100001";
Trees_din <= "00000100000000000101111100000100";
wait for Clk_period;
Addr <= "1000001100010";
Trees_din <= "00000000000111010100001001110001";
wait for Clk_period;
Addr <= "1000001100011";
Trees_din <= "00000000000010100100001001110001";
wait for Clk_period;
Addr <= "1000001100100";
Trees_din <= "00000000000000000001111100000100";
wait for Clk_period;
Addr <= "1000001100101";
Trees_din <= "00000000010101110100001001110001";
wait for Clk_period;
Addr <= "1000001100110";
Trees_din <= "00000000000111110100001001110001";
wait for Clk_period;
Addr <= "1000001100111";
Trees_din <= "00000011000000000000100100001000";
wait for Clk_period;
Addr <= "1000001101000";
Trees_din <= "00000011000000000000011100000100";
wait for Clk_period;
Addr <= "1000001101001";
Trees_din <= "00000000000101010100001001110001";
wait for Clk_period;
Addr <= "1000001101010";
Trees_din <= "00000000010101000100001001110001";
wait for Clk_period;
Addr <= "1000001101011";
Trees_din <= "00000001000000000011111000000100";
wait for Clk_period;
Addr <= "1000001101100";
Trees_din <= "00000000000100000100001001110001";
wait for Clk_period;
Addr <= "1000001101101";
Trees_din <= "00000000010010110100001001110001";
wait for Clk_period;
Addr <= "1000001101110";
Trees_din <= "00000010000000000011101000010000";
wait for Clk_period;
Addr <= "1000001101111";
Trees_din <= "00000100000000000100000000001000";
wait for Clk_period;
Addr <= "1000001110000";
Trees_din <= "00000001000000000011001100000100";
wait for Clk_period;
Addr <= "1000001110001";
Trees_din <= "00000000000011010100001001110001";
wait for Clk_period;
Addr <= "1000001110010";
Trees_din <= "00000000010101100100001001110001";
wait for Clk_period;
Addr <= "1000001110011";
Trees_din <= "00000101000000000000001000000100";
wait for Clk_period;
Addr <= "1000001110100";
Trees_din <= "00000000010101010100001001110001";
wait for Clk_period;
Addr <= "1000001110101";
Trees_din <= "00000000000110000100001001110001";
wait for Clk_period;
Addr <= "1000001110110";
Trees_din <= "00000110000000000001100000001000";
wait for Clk_period;
Addr <= "1000001110111";
Trees_din <= "00000111000000000010100000000100";
wait for Clk_period;
Addr <= "1000001111000";
Trees_din <= "00000000011000000100001001110001";
wait for Clk_period;
Addr <= "1000001111001";
Trees_din <= "00000000010111010100001001110001";
wait for Clk_period;
Addr <= "1000001111010";
Trees_din <= "00000001000000000011000000000100";
wait for Clk_period;
Addr <= "1000001111011";
Trees_din <= "00000000010001100100001001110001";
wait for Clk_period;
Addr <= "1000001111100";
Trees_din <= "00000000010100110100001001110001";
wait for Clk_period;
Addr <= "1000001111101";
Trees_din <= "00000101000000000100110000100000";
wait for Clk_period;
Addr <= "1000001111110";
Trees_din <= "00000100000000000001101100010000";
wait for Clk_period;
Addr <= "1000001111111";
Trees_din <= "00000101000000000101111100001000";
wait for Clk_period;
Addr <= "1000010000000";
Trees_din <= "00000101000000000100111100000100";
wait for Clk_period;
Addr <= "1000010000001";
Trees_din <= "00000000010010110100001001110001";
wait for Clk_period;
Addr <= "1000010000010";
Trees_din <= "00000000010011110100001001110001";
wait for Clk_period;
Addr <= "1000010000011";
Trees_din <= "00000101000000000011111100000100";
wait for Clk_period;
Addr <= "1000010000100";
Trees_din <= "00000000001100100100001001110001";
wait for Clk_period;
Addr <= "1000010000101";
Trees_din <= "00000000001111010100001001110001";
wait for Clk_period;
Addr <= "1000010000110";
Trees_din <= "00000101000000000011011100001000";
wait for Clk_period;
Addr <= "1000010000111";
Trees_din <= "00000111000000000101011100000100";
wait for Clk_period;
Addr <= "1000010001000";
Trees_din <= "00000000001100010100001001110001";
wait for Clk_period;
Addr <= "1000010001001";
Trees_din <= "00000000000100100100001001110001";
wait for Clk_period;
Addr <= "1000010001010";
Trees_din <= "00000111000000000100001000000100";
wait for Clk_period;
Addr <= "1000010001011";
Trees_din <= "00000000010110000100001001110001";
wait for Clk_period;
Addr <= "1000010001100";
Trees_din <= "00000000001101110100001001110001";
wait for Clk_period;
Addr <= "1000010001101";
Trees_din <= "00000111000000000101100000010000";
wait for Clk_period;
Addr <= "1000010001110";
Trees_din <= "00000001000000000100111100001000";
wait for Clk_period;
Addr <= "1000010001111";
Trees_din <= "00000100000000000001000000000100";
wait for Clk_period;
Addr <= "1000010010000";
Trees_din <= "00000000000000010100001001110001";
wait for Clk_period;
Addr <= "1000010010001";
Trees_din <= "00000000001011010100001001110001";
wait for Clk_period;
Addr <= "1000010010010";
Trees_din <= "00000111000000000011111000000100";
wait for Clk_period;
Addr <= "1000010010011";
Trees_din <= "00000000000001010100001001110001";
wait for Clk_period;
Addr <= "1000010010100";
Trees_din <= "00000000001000010100001001110001";
wait for Clk_period;
Addr <= "1000010010101";
Trees_din <= "00000011000000000010110000001000";
wait for Clk_period;
Addr <= "1000010010110";
Trees_din <= "00000111000000000100110000000100";
wait for Clk_period;
Addr <= "1000010010111";
Trees_din <= "00000000000101000100001001110001";
wait for Clk_period;
Addr <= "1000010011000";
Trees_din <= "00000000001111000100001001110001";
wait for Clk_period;
Addr <= "1000010011001";
Trees_din <= "00000101000000000011011100000100";
wait for Clk_period;
Addr <= "1000010011010";
Trees_din <= "00000000010001100100001001110001";
wait for Clk_period;
Addr <= "1000010011011";
Trees_din <= "00000000010001110100001001110001";
wait for Clk_period;



----------tree 33-------------------

Addr <= "1000010011100";
Trees_din <= "00000010000000000100010110000000";
wait for Clk_period;
Addr <= "1000010011101";
Trees_din <= "00000010000000000011110101000000";
wait for Clk_period;
Addr <= "1000010011110";
Trees_din <= "00000000000000000101010000100000";
wait for Clk_period;
Addr <= "1000010011111";
Trees_din <= "00000111000000000101010100010000";
wait for Clk_period;
Addr <= "1000010100000";
Trees_din <= "00000100000000000011100000001000";
wait for Clk_period;
Addr <= "1000010100001";
Trees_din <= "00000000000000000011100000000100";
wait for Clk_period;
Addr <= "1000010100010";
Trees_din <= "00000000001111000100010001101101";
wait for Clk_period;
Addr <= "1000010100011";
Trees_din <= "00000000000111100100010001101101";
wait for Clk_period;
Addr <= "1000010100100";
Trees_din <= "00000100000000000011010000000100";
wait for Clk_period;
Addr <= "1000010100101";
Trees_din <= "00000000010111000100010001101101";
wait for Clk_period;
Addr <= "1000010100110";
Trees_din <= "00000000010011110100010001101101";
wait for Clk_period;
Addr <= "1000010100111";
Trees_din <= "00000101000000000100101100001000";
wait for Clk_period;
Addr <= "1000010101000";
Trees_din <= "00000001000000000010101000000100";
wait for Clk_period;
Addr <= "1000010101001";
Trees_din <= "00000000000000100100010001101101";
wait for Clk_period;
Addr <= "1000010101010";
Trees_din <= "00000000000100110100010001101101";
wait for Clk_period;
Addr <= "1000010101011";
Trees_din <= "00000000000000000010000100000100";
wait for Clk_period;
Addr <= "1000010101100";
Trees_din <= "00000000000010010100010001101101";
wait for Clk_period;
Addr <= "1000010101101";
Trees_din <= "00000000010011000100010001101101";
wait for Clk_period;
Addr <= "1000010101110";
Trees_din <= "00000011000000000001111000010000";
wait for Clk_period;
Addr <= "1000010101111";
Trees_din <= "00000000000000000000010100001000";
wait for Clk_period;
Addr <= "1000010110000";
Trees_din <= "00000010000000000010100100000100";
wait for Clk_period;
Addr <= "1000010110001";
Trees_din <= "00000000010001110100010001101101";
wait for Clk_period;
Addr <= "1000010110010";
Trees_din <= "00000000010001000100010001101101";
wait for Clk_period;
Addr <= "1000010110011";
Trees_din <= "00000101000000000010011000000100";
wait for Clk_period;
Addr <= "1000010110100";
Trees_din <= "00000000001010010100010001101101";
wait for Clk_period;
Addr <= "1000010110101";
Trees_din <= "00000000000111010100010001101101";
wait for Clk_period;
Addr <= "1000010110110";
Trees_din <= "00000010000000000011111100001000";
wait for Clk_period;
Addr <= "1000010110111";
Trees_din <= "00000111000000000011110100000100";
wait for Clk_period;
Addr <= "1000010111000";
Trees_din <= "00000000000000110100010001101101";
wait for Clk_period;
Addr <= "1000010111001";
Trees_din <= "00000000010010010100010001101101";
wait for Clk_period;
Addr <= "1000010111010";
Trees_din <= "00000101000000000100110000000100";
wait for Clk_period;
Addr <= "1000010111011";
Trees_din <= "00000000010000100100010001101101";
wait for Clk_period;
Addr <= "1000010111100";
Trees_din <= "00000000000100000100010001101101";
wait for Clk_period;
Addr <= "1000010111101";
Trees_din <= "00000010000000000000111100100000";
wait for Clk_period;
Addr <= "1000010111110";
Trees_din <= "00000001000000000001100000010000";
wait for Clk_period;
Addr <= "1000010111111";
Trees_din <= "00000100000000000100001100001000";
wait for Clk_period;
Addr <= "1000011000000";
Trees_din <= "00000001000000000001111000000100";
wait for Clk_period;
Addr <= "1000011000001";
Trees_din <= "00000000000000010100010001101101";
wait for Clk_period;
Addr <= "1000011000010";
Trees_din <= "00000000010000010100010001101101";
wait for Clk_period;
Addr <= "1000011000011";
Trees_din <= "00000010000000000110001100000100";
wait for Clk_period;
Addr <= "1000011000100";
Trees_din <= "00000000010011110100010001101101";
wait for Clk_period;
Addr <= "1000011000101";
Trees_din <= "00000000000101010100010001101101";
wait for Clk_period;
Addr <= "1000011000110";
Trees_din <= "00000001000000000001010100001000";
wait for Clk_period;
Addr <= "1000011000111";
Trees_din <= "00000010000000000001011100000100";
wait for Clk_period;
Addr <= "1000011001000";
Trees_din <= "00000000001111110100010001101101";
wait for Clk_period;
Addr <= "1000011001001";
Trees_din <= "00000000000111100100010001101101";
wait for Clk_period;
Addr <= "1000011001010";
Trees_din <= "00000000000000000001101000000100";
wait for Clk_period;
Addr <= "1000011001011";
Trees_din <= "00000000000100000100010001101101";
wait for Clk_period;
Addr <= "1000011001100";
Trees_din <= "00000000010000010100010001101101";
wait for Clk_period;
Addr <= "1000011001101";
Trees_din <= "00000001000000000101100000010000";
wait for Clk_period;
Addr <= "1000011001110";
Trees_din <= "00000001000000000000010100001000";
wait for Clk_period;
Addr <= "1000011001111";
Trees_din <= "00000010000000000100100100000100";
wait for Clk_period;
Addr <= "1000011010000";
Trees_din <= "00000000000111110100010001101101";
wait for Clk_period;
Addr <= "1000011010001";
Trees_din <= "00000000001110010100010001101101";
wait for Clk_period;
Addr <= "1000011010010";
Trees_din <= "00000100000000000011110000000100";
wait for Clk_period;
Addr <= "1000011010011";
Trees_din <= "00000000001011000100010001101101";
wait for Clk_period;
Addr <= "1000011010100";
Trees_din <= "00000000010101110100010001101101";
wait for Clk_period;
Addr <= "1000011010101";
Trees_din <= "00000110000000000000111000001000";
wait for Clk_period;
Addr <= "1000011010110";
Trees_din <= "00000001000000000011010100000100";
wait for Clk_period;
Addr <= "1000011010111";
Trees_din <= "00000000000000100100010001101101";
wait for Clk_period;
Addr <= "1000011011000";
Trees_din <= "00000000010100010100010001101101";
wait for Clk_period;
Addr <= "1000011011001";
Trees_din <= "00000100000000000101101000000100";
wait for Clk_period;
Addr <= "1000011011010";
Trees_din <= "00000000011000110100010001101101";
wait for Clk_period;
Addr <= "1000011011011";
Trees_din <= "00000000001110110100010001101101";
wait for Clk_period;
Addr <= "1000011011100";
Trees_din <= "00000010000000000000000001000000";
wait for Clk_period;
Addr <= "1000011011101";
Trees_din <= "00000010000000000000110100100000";
wait for Clk_period;
Addr <= "1000011011110";
Trees_din <= "00000010000000000100001000010000";
wait for Clk_period;
Addr <= "1000011011111";
Trees_din <= "00000100000000000001110100001000";
wait for Clk_period;
Addr <= "1000011100000";
Trees_din <= "00000011000000000110000000000100";
wait for Clk_period;
Addr <= "1000011100001";
Trees_din <= "00000000010001000100010001101101";
wait for Clk_period;
Addr <= "1000011100010";
Trees_din <= "00000000000010110100010001101101";
wait for Clk_period;
Addr <= "1000011100011";
Trees_din <= "00000110000000000001011100000100";
wait for Clk_period;
Addr <= "1000011100100";
Trees_din <= "00000000010101010100010001101101";
wait for Clk_period;
Addr <= "1000011100101";
Trees_din <= "00000000001100100100010001101101";
wait for Clk_period;
Addr <= "1000011100110";
Trees_din <= "00000110000000000000000100001000";
wait for Clk_period;
Addr <= "1000011100111";
Trees_din <= "00000010000000000010001100000100";
wait for Clk_period;
Addr <= "1000011101000";
Trees_din <= "00000000001010000100010001101101";
wait for Clk_period;
Addr <= "1000011101001";
Trees_din <= "00000000000000100100010001101101";
wait for Clk_period;
Addr <= "1000011101010";
Trees_din <= "00000100000000000000111000000100";
wait for Clk_period;
Addr <= "1000011101011";
Trees_din <= "00000000000100010100010001101101";
wait for Clk_period;
Addr <= "1000011101100";
Trees_din <= "00000000001011110100010001101101";
wait for Clk_period;
Addr <= "1000011101101";
Trees_din <= "00000000000000000010100100010000";
wait for Clk_period;
Addr <= "1000011101110";
Trees_din <= "00000011000000000000100000001000";
wait for Clk_period;
Addr <= "1000011101111";
Trees_din <= "00000010000000000100000000000100";
wait for Clk_period;
Addr <= "1000011110000";
Trees_din <= "00000000000110010100010001101101";
wait for Clk_period;
Addr <= "1000011110001";
Trees_din <= "00000000011000100100010001101101";
wait for Clk_period;
Addr <= "1000011110010";
Trees_din <= "00000110000000000101000000000100";
wait for Clk_period;
Addr <= "1000011110011";
Trees_din <= "00000000010111100100010001101101";
wait for Clk_period;
Addr <= "1000011110100";
Trees_din <= "00000000000000110100010001101101";
wait for Clk_period;
Addr <= "1000011110101";
Trees_din <= "00000011000000000000111000001000";
wait for Clk_period;
Addr <= "1000011110110";
Trees_din <= "00000000000000000001111000000100";
wait for Clk_period;
Addr <= "1000011110111";
Trees_din <= "00000000001010000100010001101101";
wait for Clk_period;
Addr <= "1000011111000";
Trees_din <= "00000000001111000100010001101101";
wait for Clk_period;
Addr <= "1000011111001";
Trees_din <= "00000010000000000011100000000100";
wait for Clk_period;
Addr <= "1000011111010";
Trees_din <= "00000000000001100100010001101101";
wait for Clk_period;
Addr <= "1000011111011";
Trees_din <= "00000000000101010100010001101101";
wait for Clk_period;
Addr <= "1000011111100";
Trees_din <= "00000110000000000101110100100000";
wait for Clk_period;
Addr <= "1000011111101";
Trees_din <= "00000000000000000100010000010000";
wait for Clk_period;
Addr <= "1000011111110";
Trees_din <= "00000100000000000000011000001000";
wait for Clk_period;
Addr <= "1000011111111";
Trees_din <= "00000000000000000011011000000100";
wait for Clk_period;
Addr <= "1000100000000";
Trees_din <= "00000000010001000100010001101101";
wait for Clk_period;
Addr <= "1000100000001";
Trees_din <= "00000000001010100100010001101101";
wait for Clk_period;
Addr <= "1000100000010";
Trees_din <= "00000101000000000011100100000100";
wait for Clk_period;
Addr <= "1000100000011";
Trees_din <= "00000000000001000100010001101101";
wait for Clk_period;
Addr <= "1000100000100";
Trees_din <= "00000000000001110100010001101101";
wait for Clk_period;
Addr <= "1000100000101";
Trees_din <= "00000010000000000110001100001000";
wait for Clk_period;
Addr <= "1000100000110";
Trees_din <= "00000101000000000001000000000100";
wait for Clk_period;
Addr <= "1000100000111";
Trees_din <= "00000000011000100100010001101101";
wait for Clk_period;
Addr <= "1000100001000";
Trees_din <= "00000000000111100100010001101101";
wait for Clk_period;
Addr <= "1000100001001";
Trees_din <= "00000101000000000100111000000100";
wait for Clk_period;
Addr <= "1000100001010";
Trees_din <= "00000000000000100100010001101101";
wait for Clk_period;
Addr <= "1000100001011";
Trees_din <= "00000000001111000100010001101101";
wait for Clk_period;
Addr <= "1000100001100";
Trees_din <= "00000110000000000100111000010000";
wait for Clk_period;
Addr <= "1000100001101";
Trees_din <= "00000001000000000010100000001000";
wait for Clk_period;
Addr <= "1000100001110";
Trees_din <= "00000010000000000110001100000100";
wait for Clk_period;
Addr <= "1000100001111";
Trees_din <= "00000000000110110100010001101101";
wait for Clk_period;
Addr <= "1000100010000";
Trees_din <= "00000000011000000100010001101101";
wait for Clk_period;
Addr <= "1000100010001";
Trees_din <= "00000011000000000011100000000100";
wait for Clk_period;
Addr <= "1000100010010";
Trees_din <= "00000000000111010100010001101101";
wait for Clk_period;
Addr <= "1000100010011";
Trees_din <= "00000000010001110100010001101101";
wait for Clk_period;
Addr <= "1000100010100";
Trees_din <= "00000010000000000100100100001000";
wait for Clk_period;
Addr <= "1000100010101";
Trees_din <= "00000001000000000011010000000100";
wait for Clk_period;
Addr <= "1000100010110";
Trees_din <= "00000000010110010100010001101101";
wait for Clk_period;
Addr <= "1000100010111";
Trees_din <= "00000000000011110100010001101101";
wait for Clk_period;
Addr <= "1000100011000";
Trees_din <= "00000001000000000101100100000100";
wait for Clk_period;
Addr <= "1000100011001";
Trees_din <= "00000000010111010100010001101101";
wait for Clk_period;
Addr <= "1000100011010";
Trees_din <= "00000000010100110100010001101101";
wait for Clk_period;



----------tree 34-------------------

Addr <= "1000100011011";
Trees_din <= "00000111000000000100001010000000";
wait for Clk_period;
Addr <= "1000100011100";
Trees_din <= "00000001000000000100100101000000";
wait for Clk_period;
Addr <= "1000100011101";
Trees_din <= "00000110000000000010000100100000";
wait for Clk_period;
Addr <= "1000100011110";
Trees_din <= "00000110000000000101000100010000";
wait for Clk_period;
Addr <= "1000100011111";
Trees_din <= "00000100000000000100010100001000";
wait for Clk_period;
Addr <= "1000100100000";
Trees_din <= "00000000000000000101001000000100";
wait for Clk_period;
Addr <= "1000100100001";
Trees_din <= "00000000000000010100011001101001";
wait for Clk_period;
Addr <= "1000100100010";
Trees_din <= "00000000001001100100011001101001";
wait for Clk_period;
Addr <= "1000100100011";
Trees_din <= "00000001000000000100011000000100";
wait for Clk_period;
Addr <= "1000100100100";
Trees_din <= "00000000001010100100011001101001";
wait for Clk_period;
Addr <= "1000100100101";
Trees_din <= "00000000000011010100011001101001";
wait for Clk_period;
Addr <= "1000100100110";
Trees_din <= "00000011000000000011000100001000";
wait for Clk_period;
Addr <= "1000100100111";
Trees_din <= "00000111000000000100001100000100";
wait for Clk_period;
Addr <= "1000100101000";
Trees_din <= "00000000001111000100011001101001";
wait for Clk_period;
Addr <= "1000100101001";
Trees_din <= "00000000010001110100011001101001";
wait for Clk_period;
Addr <= "1000100101010";
Trees_din <= "00000110000000000101111000000100";
wait for Clk_period;
Addr <= "1000100101011";
Trees_din <= "00000000010011010100011001101001";
wait for Clk_period;
Addr <= "1000100101100";
Trees_din <= "00000000010101110100011001101001";
wait for Clk_period;
Addr <= "1000100101101";
Trees_din <= "00000001000000000001011100010000";
wait for Clk_period;
Addr <= "1000100101110";
Trees_din <= "00000000000000000100011100001000";
wait for Clk_period;
Addr <= "1000100101111";
Trees_din <= "00000011000000000010010100000100";
wait for Clk_period;
Addr <= "1000100110000";
Trees_din <= "00000000001111100100011001101001";
wait for Clk_period;
Addr <= "1000100110001";
Trees_din <= "00000000000110000100011001101001";
wait for Clk_period;
Addr <= "1000100110010";
Trees_din <= "00000110000000000110000000000100";
wait for Clk_period;
Addr <= "1000100110011";
Trees_din <= "00000000001010100100011001101001";
wait for Clk_period;
Addr <= "1000100110100";
Trees_din <= "00000000010011010100011001101001";
wait for Clk_period;
Addr <= "1000100110101";
Trees_din <= "00000010000000000001011100001000";
wait for Clk_period;
Addr <= "1000100110110";
Trees_din <= "00000100000000000001011100000100";
wait for Clk_period;
Addr <= "1000100110111";
Trees_din <= "00000000001010110100011001101001";
wait for Clk_period;
Addr <= "1000100111000";
Trees_din <= "00000000000010100100011001101001";
wait for Clk_period;
Addr <= "1000100111001";
Trees_din <= "00000010000000000101001100000100";
wait for Clk_period;
Addr <= "1000100111010";
Trees_din <= "00000000001100010100011001101001";
wait for Clk_period;
Addr <= "1000100111011";
Trees_din <= "00000000001011100100011001101001";
wait for Clk_period;
Addr <= "1000100111100";
Trees_din <= "00000111000000000110001000100000";
wait for Clk_period;
Addr <= "1000100111101";
Trees_din <= "00000000000000000011010000010000";
wait for Clk_period;
Addr <= "1000100111110";
Trees_din <= "00000011000000000011100100001000";
wait for Clk_period;
Addr <= "1000100111111";
Trees_din <= "00000010000000000000100100000100";
wait for Clk_period;
Addr <= "1000101000000";
Trees_din <= "00000000000101110100011001101001";
wait for Clk_period;
Addr <= "1000101000001";
Trees_din <= "00000000001011110100011001101001";
wait for Clk_period;
Addr <= "1000101000010";
Trees_din <= "00000010000000000001001000000100";
wait for Clk_period;
Addr <= "1000101000011";
Trees_din <= "00000000000001010100011001101001";
wait for Clk_period;
Addr <= "1000101000100";
Trees_din <= "00000000010010010100011001101001";
wait for Clk_period;
Addr <= "1000101000101";
Trees_din <= "00000101000000000101001000001000";
wait for Clk_period;
Addr <= "1000101000110";
Trees_din <= "00000101000000000001110100000100";
wait for Clk_period;
Addr <= "1000101000111";
Trees_din <= "00000000001010010100011001101001";
wait for Clk_period;
Addr <= "1000101001000";
Trees_din <= "00000000000110010100011001101001";
wait for Clk_period;
Addr <= "1000101001001";
Trees_din <= "00000101000000000000110100000100";
wait for Clk_period;
Addr <= "1000101001010";
Trees_din <= "00000000010110100100011001101001";
wait for Clk_period;
Addr <= "1000101001011";
Trees_din <= "00000000001000010100011001101001";
wait for Clk_period;
Addr <= "1000101001100";
Trees_din <= "00000101000000000101101000010000";
wait for Clk_period;
Addr <= "1000101001101";
Trees_din <= "00000100000000000001001000001000";
wait for Clk_period;
Addr <= "1000101001110";
Trees_din <= "00000101000000000001010100000100";
wait for Clk_period;
Addr <= "1000101001111";
Trees_din <= "00000000000100010100011001101001";
wait for Clk_period;
Addr <= "1000101010000";
Trees_din <= "00000000010011010100011001101001";
wait for Clk_period;
Addr <= "1000101010001";
Trees_din <= "00000011000000000100001100000100";
wait for Clk_period;
Addr <= "1000101010010";
Trees_din <= "00000000001011110100011001101001";
wait for Clk_period;
Addr <= "1000101010011";
Trees_din <= "00000000010011000100011001101001";
wait for Clk_period;
Addr <= "1000101010100";
Trees_din <= "00000101000000000011101000001000";
wait for Clk_period;
Addr <= "1000101010101";
Trees_din <= "00000010000000000010110000000100";
wait for Clk_period;
Addr <= "1000101010110";
Trees_din <= "00000000010000110100011001101001";
wait for Clk_period;
Addr <= "1000101010111";
Trees_din <= "00000000001001010100011001101001";
wait for Clk_period;
Addr <= "1000101011000";
Trees_din <= "00000000000000000010000100000100";
wait for Clk_period;
Addr <= "1000101011001";
Trees_din <= "00000000001110100100011001101001";
wait for Clk_period;
Addr <= "1000101011010";
Trees_din <= "00000000010101010100011001101001";
wait for Clk_period;
Addr <= "1000101011011";
Trees_din <= "00000000000000000001111101000000";
wait for Clk_period;
Addr <= "1000101011100";
Trees_din <= "00000110000000000110010000100000";
wait for Clk_period;
Addr <= "1000101011101";
Trees_din <= "00000100000000000100110000010000";
wait for Clk_period;
Addr <= "1000101011110";
Trees_din <= "00000001000000000010001100001000";
wait for Clk_period;
Addr <= "1000101011111";
Trees_din <= "00000000000000000000001100000100";
wait for Clk_period;
Addr <= "1000101100000";
Trees_din <= "00000000000100110100011001101001";
wait for Clk_period;
Addr <= "1000101100001";
Trees_din <= "00000000001110100100011001101001";
wait for Clk_period;
Addr <= "1000101100010";
Trees_din <= "00000111000000000001010100000100";
wait for Clk_period;
Addr <= "1000101100011";
Trees_din <= "00000000000110100100011001101001";
wait for Clk_period;
Addr <= "1000101100100";
Trees_din <= "00000000000110110100011001101001";
wait for Clk_period;
Addr <= "1000101100101";
Trees_din <= "00000000000000000101101100001000";
wait for Clk_period;
Addr <= "1000101100110";
Trees_din <= "00000101000000000001110100000100";
wait for Clk_period;
Addr <= "1000101100111";
Trees_din <= "00000000011000010100011001101001";
wait for Clk_period;
Addr <= "1000101101000";
Trees_din <= "00000000010110100100011001101001";
wait for Clk_period;
Addr <= "1000101101001";
Trees_din <= "00000010000000000011110100000100";
wait for Clk_period;
Addr <= "1000101101010";
Trees_din <= "00000000010001000100011001101001";
wait for Clk_period;
Addr <= "1000101101011";
Trees_din <= "00000000010101110100011001101001";
wait for Clk_period;
Addr <= "1000101101100";
Trees_din <= "00000011000000000100100100010000";
wait for Clk_period;
Addr <= "1000101101101";
Trees_din <= "00000101000000000010001100001000";
wait for Clk_period;
Addr <= "1000101101110";
Trees_din <= "00000011000000000101110100000100";
wait for Clk_period;
Addr <= "1000101101111";
Trees_din <= "00000000010011010100011001101001";
wait for Clk_period;
Addr <= "1000101110000";
Trees_din <= "00000000011000110100011001101001";
wait for Clk_period;
Addr <= "1000101110001";
Trees_din <= "00000000000000000000011100000100";
wait for Clk_period;
Addr <= "1000101110010";
Trees_din <= "00000000000110010100011001101001";
wait for Clk_period;
Addr <= "1000101110011";
Trees_din <= "00000000001000010100011001101001";
wait for Clk_period;
Addr <= "1000101110100";
Trees_din <= "00000000000000000011011100001000";
wait for Clk_period;
Addr <= "1000101110101";
Trees_din <= "00000001000000000000111000000100";
wait for Clk_period;
Addr <= "1000101110110";
Trees_din <= "00000000001011100100011001101001";
wait for Clk_period;
Addr <= "1000101110111";
Trees_din <= "00000000000110000100011001101001";
wait for Clk_period;
Addr <= "1000101111000";
Trees_din <= "00000110000000000010001000000100";
wait for Clk_period;
Addr <= "1000101111001";
Trees_din <= "00000000000101010100011001101001";
wait for Clk_period;
Addr <= "1000101111010";
Trees_din <= "00000000001111100100011001101001";
wait for Clk_period;
Addr <= "1000101111011";
Trees_din <= "00000100000000000001110100100000";
wait for Clk_period;
Addr <= "1000101111100";
Trees_din <= "00000101000000000100101000010000";
wait for Clk_period;
Addr <= "1000101111101";
Trees_din <= "00000000000000000000001000001000";
wait for Clk_period;
Addr <= "1000101111110";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "1000101111111";
Trees_din <= "00000000001111100100011001101001";
wait for Clk_period;
Addr <= "1000110000000";
Trees_din <= "00000000010100000100011001101001";
wait for Clk_period;
Addr <= "1000110000001";
Trees_din <= "00000001000000000001000100000100";
wait for Clk_period;
Addr <= "1000110000010";
Trees_din <= "00000000010100110100011001101001";
wait for Clk_period;
Addr <= "1000110000011";
Trees_din <= "00000000001111010100011001101001";
wait for Clk_period;
Addr <= "1000110000100";
Trees_din <= "00000011000000000000101000001000";
wait for Clk_period;
Addr <= "1000110000101";
Trees_din <= "00000011000000000000111100000100";
wait for Clk_period;
Addr <= "1000110000110";
Trees_din <= "00000000001011110100011001101001";
wait for Clk_period;
Addr <= "1000110000111";
Trees_din <= "00000000011000010100011001101001";
wait for Clk_period;
Addr <= "1000110001000";
Trees_din <= "00000101000000000000001000000100";
wait for Clk_period;
Addr <= "1000110001001";
Trees_din <= "00000000010101010100011001101001";
wait for Clk_period;
Addr <= "1000110001010";
Trees_din <= "00000000001111100100011001101001";
wait for Clk_period;
Addr <= "1000110001011";
Trees_din <= "00000110000000000101000000010000";
wait for Clk_period;
Addr <= "1000110001100";
Trees_din <= "00000101000000000000100100001000";
wait for Clk_period;
Addr <= "1000110001101";
Trees_din <= "00000111000000000011101000000100";
wait for Clk_period;
Addr <= "1000110001110";
Trees_din <= "00000000010011110100011001101001";
wait for Clk_period;
Addr <= "1000110001111";
Trees_din <= "00000000001000100100011001101001";
wait for Clk_period;
Addr <= "1000110010000";
Trees_din <= "00000000000000000011101100000100";
wait for Clk_period;
Addr <= "1000110010001";
Trees_din <= "00000000001111000100011001101001";
wait for Clk_period;
Addr <= "1000110010010";
Trees_din <= "00000000001110110100011001101001";
wait for Clk_period;
Addr <= "1000110010011";
Trees_din <= "00000011000000000100010100001000";
wait for Clk_period;
Addr <= "1000110010100";
Trees_din <= "00000000000000000010110100000100";
wait for Clk_period;
Addr <= "1000110010101";
Trees_din <= "00000000000100000100011001101001";
wait for Clk_period;
Addr <= "1000110010110";
Trees_din <= "00000000001000110100011001101001";
wait for Clk_period;
Addr <= "1000110010111";
Trees_din <= "00000010000000000011011000000100";
wait for Clk_period;
Addr <= "1000110011000";
Trees_din <= "00000000010001110100011001101001";
wait for Clk_period;
Addr <= "1000110011001";
Trees_din <= "00000000001110010100011001101001";
wait for Clk_period;



----------tree 35-------------------

Addr <= "1000110011010";
Trees_din <= "00000100000000000011101110000000";
wait for Clk_period;
Addr <= "1000110011011";
Trees_din <= "00000111000000000001111001000000";
wait for Clk_period;
Addr <= "1000110011100";
Trees_din <= "00000100000000000001001000100000";
wait for Clk_period;
Addr <= "1000110011101";
Trees_din <= "00000001000000000011101000010000";
wait for Clk_period;
Addr <= "1000110011110";
Trees_din <= "00000011000000000011001100001000";
wait for Clk_period;
Addr <= "1000110011111";
Trees_din <= "00000010000000000011010100000100";
wait for Clk_period;
Addr <= "1000110100000";
Trees_din <= "00000000011000000100100001100101";
wait for Clk_period;
Addr <= "1000110100001";
Trees_din <= "00000000010110100100100001100101";
wait for Clk_period;
Addr <= "1000110100010";
Trees_din <= "00000101000000000011010000000100";
wait for Clk_period;
Addr <= "1000110100011";
Trees_din <= "00000000001001100100100001100101";
wait for Clk_period;
Addr <= "1000110100100";
Trees_din <= "00000000010001100100100001100101";
wait for Clk_period;
Addr <= "1000110100101";
Trees_din <= "00000000000000000001001000001000";
wait for Clk_period;
Addr <= "1000110100110";
Trees_din <= "00000000000000000000001100000100";
wait for Clk_period;
Addr <= "1000110100111";
Trees_din <= "00000000011000110100100001100101";
wait for Clk_period;
Addr <= "1000110101000";
Trees_din <= "00000000001101100100100001100101";
wait for Clk_period;
Addr <= "1000110101001";
Trees_din <= "00000001000000000100111100000100";
wait for Clk_period;
Addr <= "1000110101010";
Trees_din <= "00000000001011110100100001100101";
wait for Clk_period;
Addr <= "1000110101011";
Trees_din <= "00000000000111100100100001100101";
wait for Clk_period;
Addr <= "1000110101100";
Trees_din <= "00000111000000000100101000010000";
wait for Clk_period;
Addr <= "1000110101101";
Trees_din <= "00000110000000000001110100001000";
wait for Clk_period;
Addr <= "1000110101110";
Trees_din <= "00000011000000000000010100000100";
wait for Clk_period;
Addr <= "1000110101111";
Trees_din <= "00000000001001000100100001100101";
wait for Clk_period;
Addr <= "1000110110000";
Trees_din <= "00000000000100100100100001100101";
wait for Clk_period;
Addr <= "1000110110001";
Trees_din <= "00000111000000000100010000000100";
wait for Clk_period;
Addr <= "1000110110010";
Trees_din <= "00000000000111010100100001100101";
wait for Clk_period;
Addr <= "1000110110011";
Trees_din <= "00000000010011000100100001100101";
wait for Clk_period;
Addr <= "1000110110100";
Trees_din <= "00000111000000000011111100001000";
wait for Clk_period;
Addr <= "1000110110101";
Trees_din <= "00000010000000000101111100000100";
wait for Clk_period;
Addr <= "1000110110110";
Trees_din <= "00000000011000100100100001100101";
wait for Clk_period;
Addr <= "1000110110111";
Trees_din <= "00000000011000000100100001100101";
wait for Clk_period;
Addr <= "1000110111000";
Trees_din <= "00000100000000000010111000000100";
wait for Clk_period;
Addr <= "1000110111001";
Trees_din <= "00000000000010010100100001100101";
wait for Clk_period;
Addr <= "1000110111010";
Trees_din <= "00000000001110110100100001100101";
wait for Clk_period;
Addr <= "1000110111011";
Trees_din <= "00000111000000000100101100100000";
wait for Clk_period;
Addr <= "1000110111100";
Trees_din <= "00000101000000000010101000010000";
wait for Clk_period;
Addr <= "1000110111101";
Trees_din <= "00000100000000000110001000001000";
wait for Clk_period;
Addr <= "1000110111110";
Trees_din <= "00000001000000000011001000000100";
wait for Clk_period;
Addr <= "1000110111111";
Trees_din <= "00000000010110110100100001100101";
wait for Clk_period;
Addr <= "1000111000000";
Trees_din <= "00000000001100100100100001100101";
wait for Clk_period;
Addr <= "1000111000001";
Trees_din <= "00000111000000000100100100000100";
wait for Clk_period;
Addr <= "1000111000010";
Trees_din <= "00000000000000110100100001100101";
wait for Clk_period;
Addr <= "1000111000011";
Trees_din <= "00000000010001100100100001100101";
wait for Clk_period;
Addr <= "1000111000100";
Trees_din <= "00000110000000000001100100001000";
wait for Clk_period;
Addr <= "1000111000101";
Trees_din <= "00000101000000000010010100000100";
wait for Clk_period;
Addr <= "1000111000110";
Trees_din <= "00000000001010000100100001100101";
wait for Clk_period;
Addr <= "1000111000111";
Trees_din <= "00000000000000110100100001100101";
wait for Clk_period;
Addr <= "1000111001000";
Trees_din <= "00000000000000000001011100000100";
wait for Clk_period;
Addr <= "1000111001001";
Trees_din <= "00000000001101110100100001100101";
wait for Clk_period;
Addr <= "1000111001010";
Trees_din <= "00000000000111010100100001100101";
wait for Clk_period;
Addr <= "1000111001011";
Trees_din <= "00000001000000000001001000010000";
wait for Clk_period;
Addr <= "1000111001100";
Trees_din <= "00000010000000000001111000001000";
wait for Clk_period;
Addr <= "1000111001101";
Trees_din <= "00000110000000000010101000000100";
wait for Clk_period;
Addr <= "1000111001110";
Trees_din <= "00000000000000010100100001100101";
wait for Clk_period;
Addr <= "1000111001111";
Trees_din <= "00000000010000110100100001100101";
wait for Clk_period;
Addr <= "1000111010000";
Trees_din <= "00000010000000000010101000000100";
wait for Clk_period;
Addr <= "1000111010001";
Trees_din <= "00000000000010000100100001100101";
wait for Clk_period;
Addr <= "1000111010010";
Trees_din <= "00000000001101110100100001100101";
wait for Clk_period;
Addr <= "1000111010011";
Trees_din <= "00000010000000000011000000001000";
wait for Clk_period;
Addr <= "1000111010100";
Trees_din <= "00000011000000000010100000000100";
wait for Clk_period;
Addr <= "1000111010101";
Trees_din <= "00000000001011110100100001100101";
wait for Clk_period;
Addr <= "1000111010110";
Trees_din <= "00000000000011110100100001100101";
wait for Clk_period;
Addr <= "1000111010111";
Trees_din <= "00000010000000000100111000000100";
wait for Clk_period;
Addr <= "1000111011000";
Trees_din <= "00000000001010100100100001100101";
wait for Clk_period;
Addr <= "1000111011001";
Trees_din <= "00000000010101010100100001100101";
wait for Clk_period;
Addr <= "1000111011010";
Trees_din <= "00000110000000000000101001000000";
wait for Clk_period;
Addr <= "1000111011011";
Trees_din <= "00000110000000000011000000100000";
wait for Clk_period;
Addr <= "1000111011100";
Trees_din <= "00000010000000000110000000010000";
wait for Clk_period;
Addr <= "1000111011101";
Trees_din <= "00000110000000000011100100001000";
wait for Clk_period;
Addr <= "1000111011110";
Trees_din <= "00000111000000000001101000000100";
wait for Clk_period;
Addr <= "1000111011111";
Trees_din <= "00000000001101100100100001100101";
wait for Clk_period;
Addr <= "1000111100000";
Trees_din <= "00000000000000000100100001100101";
wait for Clk_period;
Addr <= "1000111100001";
Trees_din <= "00000010000000000010001000000100";
wait for Clk_period;
Addr <= "1000111100010";
Trees_din <= "00000000000111000100100001100101";
wait for Clk_period;
Addr <= "1000111100011";
Trees_din <= "00000000000001100100100001100101";
wait for Clk_period;
Addr <= "1000111100100";
Trees_din <= "00000100000000000100110100001000";
wait for Clk_period;
Addr <= "1000111100101";
Trees_din <= "00000001000000000101111000000100";
wait for Clk_period;
Addr <= "1000111100110";
Trees_din <= "00000000011000110100100001100101";
wait for Clk_period;
Addr <= "1000111100111";
Trees_din <= "00000000001010110100100001100101";
wait for Clk_period;
Addr <= "1000111101000";
Trees_din <= "00000010000000000000111000000100";
wait for Clk_period;
Addr <= "1000111101001";
Trees_din <= "00000000001001000100100001100101";
wait for Clk_period;
Addr <= "1000111101010";
Trees_din <= "00000000000000010100100001100101";
wait for Clk_period;
Addr <= "1000111101011";
Trees_din <= "00000101000000000100000000010000";
wait for Clk_period;
Addr <= "1000111101100";
Trees_din <= "00000101000000000000001000001000";
wait for Clk_period;
Addr <= "1000111101101";
Trees_din <= "00000010000000000101101000000100";
wait for Clk_period;
Addr <= "1000111101110";
Trees_din <= "00000000000001000100100001100101";
wait for Clk_period;
Addr <= "1000111101111";
Trees_din <= "00000000010110110100100001100101";
wait for Clk_period;
Addr <= "1000111110000";
Trees_din <= "00000011000000000000110100000100";
wait for Clk_period;
Addr <= "1000111110001";
Trees_din <= "00000000010010110100100001100101";
wait for Clk_period;
Addr <= "1000111110010";
Trees_din <= "00000000000111010100100001100101";
wait for Clk_period;
Addr <= "1000111110011";
Trees_din <= "00000110000000000011000100001000";
wait for Clk_period;
Addr <= "1000111110100";
Trees_din <= "00000111000000000010001000000100";
wait for Clk_period;
Addr <= "1000111110101";
Trees_din <= "00000000000010010100100001100101";
wait for Clk_period;
Addr <= "1000111110110";
Trees_din <= "00000000010110100100100001100101";
wait for Clk_period;
Addr <= "1000111110111";
Trees_din <= "00000101000000000101000100000100";
wait for Clk_period;
Addr <= "1000111111000";
Trees_din <= "00000000001000000100100001100101";
wait for Clk_period;
Addr <= "1000111111001";
Trees_din <= "00000000010001100100100001100101";
wait for Clk_period;
Addr <= "1000111111010";
Trees_din <= "00000011000000000101001000100000";
wait for Clk_period;
Addr <= "1000111111011";
Trees_din <= "00000011000000000100001100010000";
wait for Clk_period;
Addr <= "1000111111100";
Trees_din <= "00000111000000000010010000001000";
wait for Clk_period;
Addr <= "1000111111101";
Trees_din <= "00000000000000000100100000000100";
wait for Clk_period;
Addr <= "1000111111110";
Trees_din <= "00000000000010010100100001100101";
wait for Clk_period;
Addr <= "1000111111111";
Trees_din <= "00000000001001010100100001100101";
wait for Clk_period;
Addr <= "1001000000000";
Trees_din <= "00000110000000000011110100000100";
wait for Clk_period;
Addr <= "1001000000001";
Trees_din <= "00000000000001000100100001100101";
wait for Clk_period;
Addr <= "1001000000010";
Trees_din <= "00000000001111100100100001100101";
wait for Clk_period;
Addr <= "1001000000011";
Trees_din <= "00000010000000000001110100001000";
wait for Clk_period;
Addr <= "1001000000100";
Trees_din <= "00000111000000000000101000000100";
wait for Clk_period;
Addr <= "1001000000101";
Trees_din <= "00000000000011010100100001100101";
wait for Clk_period;
Addr <= "1001000000110";
Trees_din <= "00000000000000110100100001100101";
wait for Clk_period;
Addr <= "1001000000111";
Trees_din <= "00000001000000000001011000000100";
wait for Clk_period;
Addr <= "1001000001000";
Trees_din <= "00000000001100000100100001100101";
wait for Clk_period;
Addr <= "1001000001001";
Trees_din <= "00000000001010100100100001100101";
wait for Clk_period;
Addr <= "1001000001010";
Trees_din <= "00000010000000000001101100010000";
wait for Clk_period;
Addr <= "1001000001011";
Trees_din <= "00000111000000000101011000001000";
wait for Clk_period;
Addr <= "1001000001100";
Trees_din <= "00000111000000000000010100000100";
wait for Clk_period;
Addr <= "1001000001101";
Trees_din <= "00000000001111000100100001100101";
wait for Clk_period;
Addr <= "1001000001110";
Trees_din <= "00000000001111100100100001100101";
wait for Clk_period;
Addr <= "1001000001111";
Trees_din <= "00000010000000000100010000000100";
wait for Clk_period;
Addr <= "1001000010000";
Trees_din <= "00000000000010000100100001100101";
wait for Clk_period;
Addr <= "1001000010001";
Trees_din <= "00000000000010000100100001100101";
wait for Clk_period;
Addr <= "1001000010010";
Trees_din <= "00000001000000000011110000001000";
wait for Clk_period;
Addr <= "1001000010011";
Trees_din <= "00000011000000000010110100000100";
wait for Clk_period;
Addr <= "1001000010100";
Trees_din <= "00000000000010110100100001100101";
wait for Clk_period;
Addr <= "1001000010101";
Trees_din <= "00000000001111010100100001100101";
wait for Clk_period;
Addr <= "1001000010110";
Trees_din <= "00000010000000000001101100000100";
wait for Clk_period;
Addr <= "1001000010111";
Trees_din <= "00000000010110100100100001100101";
wait for Clk_period;
Addr <= "1001000011000";
Trees_din <= "00000000001110100100100001100101";
wait for Clk_period;



----------tree 36-------------------

Addr <= "1001000011001";
Trees_din <= "00000000000000000101001110000000";
wait for Clk_period;
Addr <= "1001000011010";
Trees_din <= "00000011000000000011110101000000";
wait for Clk_period;
Addr <= "1001000011011";
Trees_din <= "00000110000000000000011000100000";
wait for Clk_period;
Addr <= "1001000011100";
Trees_din <= "00000011000000000010110000010000";
wait for Clk_period;
Addr <= "1001000011101";
Trees_din <= "00000111000000000100010100001000";
wait for Clk_period;
Addr <= "1001000011110";
Trees_din <= "00000100000000000011111000000100";
wait for Clk_period;
Addr <= "1001000011111";
Trees_din <= "00000000010101100100101001100001";
wait for Clk_period;
Addr <= "1001000100000";
Trees_din <= "00000000001110110100101001100001";
wait for Clk_period;
Addr <= "1001000100001";
Trees_din <= "00000001000000000010101100000100";
wait for Clk_period;
Addr <= "1001000100010";
Trees_din <= "00000000001010110100101001100001";
wait for Clk_period;
Addr <= "1001000100011";
Trees_din <= "00000000010110000100101001100001";
wait for Clk_period;
Addr <= "1001000100100";
Trees_din <= "00000110000000000110000000001000";
wait for Clk_period;
Addr <= "1001000100101";
Trees_din <= "00000101000000000001011000000100";
wait for Clk_period;
Addr <= "1001000100110";
Trees_din <= "00000000001101110100101001100001";
wait for Clk_period;
Addr <= "1001000100111";
Trees_din <= "00000000010000100100101001100001";
wait for Clk_period;
Addr <= "1001000101000";
Trees_din <= "00000101000000000101101000000100";
wait for Clk_period;
Addr <= "1001000101001";
Trees_din <= "00000000000011010100101001100001";
wait for Clk_period;
Addr <= "1001000101010";
Trees_din <= "00000000000010110100101001100001";
wait for Clk_period;
Addr <= "1001000101011";
Trees_din <= "00000010000000000000001100010000";
wait for Clk_period;
Addr <= "1001000101100";
Trees_din <= "00000111000000000010100100001000";
wait for Clk_period;
Addr <= "1001000101101";
Trees_din <= "00000010000000000100001000000100";
wait for Clk_period;
Addr <= "1001000101110";
Trees_din <= "00000000001101110100101001100001";
wait for Clk_period;
Addr <= "1001000101111";
Trees_din <= "00000000001101100100101001100001";
wait for Clk_period;
Addr <= "1001000110000";
Trees_din <= "00000100000000000100101000000100";
wait for Clk_period;
Addr <= "1001000110001";
Trees_din <= "00000000011001000100101001100001";
wait for Clk_period;
Addr <= "1001000110010";
Trees_din <= "00000000001100110100101001100001";
wait for Clk_period;
Addr <= "1001000110011";
Trees_din <= "00000100000000000100111000001000";
wait for Clk_period;
Addr <= "1001000110100";
Trees_din <= "00000001000000000011011100000100";
wait for Clk_period;
Addr <= "1001000110101";
Trees_din <= "00000000010110010100101001100001";
wait for Clk_period;
Addr <= "1001000110110";
Trees_din <= "00000000001111000100101001100001";
wait for Clk_period;
Addr <= "1001000110111";
Trees_din <= "00000111000000000001110000000100";
wait for Clk_period;
Addr <= "1001000111000";
Trees_din <= "00000000011001000100101001100001";
wait for Clk_period;
Addr <= "1001000111001";
Trees_din <= "00000000010101000100101001100001";
wait for Clk_period;
Addr <= "1001000111010";
Trees_din <= "00000111000000000101000000100000";
wait for Clk_period;
Addr <= "1001000111011";
Trees_din <= "00000111000000000001001100010000";
wait for Clk_period;
Addr <= "1001000111100";
Trees_din <= "00000100000000000101101100001000";
wait for Clk_period;
Addr <= "1001000111101";
Trees_din <= "00000111000000000000111100000100";
wait for Clk_period;
Addr <= "1001000111110";
Trees_din <= "00000000000001100100101001100001";
wait for Clk_period;
Addr <= "1001000111111";
Trees_din <= "00000000001011110100101001100001";
wait for Clk_period;
Addr <= "1001001000000";
Trees_din <= "00000000000000000000110100000100";
wait for Clk_period;
Addr <= "1001001000001";
Trees_din <= "00000000000010110100101001100001";
wait for Clk_period;
Addr <= "1001001000010";
Trees_din <= "00000000000000010100101001100001";
wait for Clk_period;
Addr <= "1001001000011";
Trees_din <= "00000000000000000010110000001000";
wait for Clk_period;
Addr <= "1001001000100";
Trees_din <= "00000111000000000000100100000100";
wait for Clk_period;
Addr <= "1001001000101";
Trees_din <= "00000000001101110100101001100001";
wait for Clk_period;
Addr <= "1001001000110";
Trees_din <= "00000000001010010100101001100001";
wait for Clk_period;
Addr <= "1001001000111";
Trees_din <= "00000101000000000100110100000100";
wait for Clk_period;
Addr <= "1001001001000";
Trees_din <= "00000000000111110100101001100001";
wait for Clk_period;
Addr <= "1001001001001";
Trees_din <= "00000000010101010100101001100001";
wait for Clk_period;
Addr <= "1001001001010";
Trees_din <= "00000100000000000100000100010000";
wait for Clk_period;
Addr <= "1001001001011";
Trees_din <= "00000011000000000000111100001000";
wait for Clk_period;
Addr <= "1001001001100";
Trees_din <= "00000001000000000101100000000100";
wait for Clk_period;
Addr <= "1001001001101";
Trees_din <= "00000000010111000100101001100001";
wait for Clk_period;
Addr <= "1001001001110";
Trees_din <= "00000000001101110100101001100001";
wait for Clk_period;
Addr <= "1001001001111";
Trees_din <= "00000111000000000100111000000100";
wait for Clk_period;
Addr <= "1001001010000";
Trees_din <= "00000000000100010100101001100001";
wait for Clk_period;
Addr <= "1001001010001";
Trees_din <= "00000000001001110100101001100001";
wait for Clk_period;
Addr <= "1001001010010";
Trees_din <= "00000001000000000101100000001000";
wait for Clk_period;
Addr <= "1001001010011";
Trees_din <= "00000010000000000100101100000100";
wait for Clk_period;
Addr <= "1001001010100";
Trees_din <= "00000000000101100100101001100001";
wait for Clk_period;
Addr <= "1001001010101";
Trees_din <= "00000000000100010100101001100001";
wait for Clk_period;
Addr <= "1001001010110";
Trees_din <= "00000111000000000101111100000100";
wait for Clk_period;
Addr <= "1001001010111";
Trees_din <= "00000000000111010100101001100001";
wait for Clk_period;
Addr <= "1001001011000";
Trees_din <= "00000000001001010100101001100001";
wait for Clk_period;
Addr <= "1001001011001";
Trees_din <= "00000011000000000011001001000000";
wait for Clk_period;
Addr <= "1001001011010";
Trees_din <= "00000111000000000110010000100000";
wait for Clk_period;
Addr <= "1001001011011";
Trees_din <= "00000101000000000001011000010000";
wait for Clk_period;
Addr <= "1001001011100";
Trees_din <= "00000011000000000110000000001000";
wait for Clk_period;
Addr <= "1001001011101";
Trees_din <= "00000001000000000000011000000100";
wait for Clk_period;
Addr <= "1001001011110";
Trees_din <= "00000000000000010100101001100001";
wait for Clk_period;
Addr <= "1001001011111";
Trees_din <= "00000000010100110100101001100001";
wait for Clk_period;
Addr <= "1001001100000";
Trees_din <= "00000101000000000010110100000100";
wait for Clk_period;
Addr <= "1001001100001";
Trees_din <= "00000000010111100100101001100001";
wait for Clk_period;
Addr <= "1001001100010";
Trees_din <= "00000000001110010100101001100001";
wait for Clk_period;
Addr <= "1001001100011";
Trees_din <= "00000110000000000011100000001000";
wait for Clk_period;
Addr <= "1001001100100";
Trees_din <= "00000110000000000000110100000100";
wait for Clk_period;
Addr <= "1001001100101";
Trees_din <= "00000000001110000100101001100001";
wait for Clk_period;
Addr <= "1001001100110";
Trees_din <= "00000000001011100100101001100001";
wait for Clk_period;
Addr <= "1001001100111";
Trees_din <= "00000111000000000000001100000100";
wait for Clk_period;
Addr <= "1001001101000";
Trees_din <= "00000000000001010100101001100001";
wait for Clk_period;
Addr <= "1001001101001";
Trees_din <= "00000000001110100100101001100001";
wait for Clk_period;
Addr <= "1001001101010";
Trees_din <= "00000001000000000101100000010000";
wait for Clk_period;
Addr <= "1001001101011";
Trees_din <= "00000110000000000010101000001000";
wait for Clk_period;
Addr <= "1001001101100";
Trees_din <= "00000011000000000011001100000100";
wait for Clk_period;
Addr <= "1001001101101";
Trees_din <= "00000000000001000100101001100001";
wait for Clk_period;
Addr <= "1001001101110";
Trees_din <= "00000000001011010100101001100001";
wait for Clk_period;
Addr <= "1001001101111";
Trees_din <= "00000100000000000000000100000100";
wait for Clk_period;
Addr <= "1001001110000";
Trees_din <= "00000000001101000100101001100001";
wait for Clk_period;
Addr <= "1001001110001";
Trees_din <= "00000000010110110100101001100001";
wait for Clk_period;
Addr <= "1001001110010";
Trees_din <= "00000111000000000101000000001000";
wait for Clk_period;
Addr <= "1001001110011";
Trees_din <= "00000110000000000100011100000100";
wait for Clk_period;
Addr <= "1001001110100";
Trees_din <= "00000000001110000100101001100001";
wait for Clk_period;
Addr <= "1001001110101";
Trees_din <= "00000000000000000100101001100001";
wait for Clk_period;
Addr <= "1001001110110";
Trees_din <= "00000111000000000100110000000100";
wait for Clk_period;
Addr <= "1001001110111";
Trees_din <= "00000000001011110100101001100001";
wait for Clk_period;
Addr <= "1001001111000";
Trees_din <= "00000000000001000100101001100001";
wait for Clk_period;
Addr <= "1001001111001";
Trees_din <= "00000000000000000000000100100000";
wait for Clk_period;
Addr <= "1001001111010";
Trees_din <= "00000011000000000000011100010000";
wait for Clk_period;
Addr <= "1001001111011";
Trees_din <= "00000100000000000001001000001000";
wait for Clk_period;
Addr <= "1001001111100";
Trees_din <= "00000111000000000000100100000100";
wait for Clk_period;
Addr <= "1001001111101";
Trees_din <= "00000000000000100100101001100001";
wait for Clk_period;
Addr <= "1001001111110";
Trees_din <= "00000000000011000100101001100001";
wait for Clk_period;
Addr <= "1001001111111";
Trees_din <= "00000110000000000000111000000100";
wait for Clk_period;
Addr <= "1001010000000";
Trees_din <= "00000000001100110100101001100001";
wait for Clk_period;
Addr <= "1001010000001";
Trees_din <= "00000000001101000100101001100001";
wait for Clk_period;
Addr <= "1001010000010";
Trees_din <= "00000011000000000011001100001000";
wait for Clk_period;
Addr <= "1001010000011";
Trees_din <= "00000000000000000010010100000100";
wait for Clk_period;
Addr <= "1001010000100";
Trees_din <= "00000000001001000100101001100001";
wait for Clk_period;
Addr <= "1001010000101";
Trees_din <= "00000000000001000100101001100001";
wait for Clk_period;
Addr <= "1001010000110";
Trees_din <= "00000000000000000100000000000100";
wait for Clk_period;
Addr <= "1001010000111";
Trees_din <= "00000000010101100100101001100001";
wait for Clk_period;
Addr <= "1001010001000";
Trees_din <= "00000000001101000100101001100001";
wait for Clk_period;
Addr <= "1001010001001";
Trees_din <= "00000110000000000100101000010000";
wait for Clk_period;
Addr <= "1001010001010";
Trees_din <= "00000100000000000110001100001000";
wait for Clk_period;
Addr <= "1001010001011";
Trees_din <= "00000000000000000100011000000100";
wait for Clk_period;
Addr <= "1001010001100";
Trees_din <= "00000000010001010100101001100001";
wait for Clk_period;
Addr <= "1001010001101";
Trees_din <= "00000000010101100100101001100001";
wait for Clk_period;
Addr <= "1001010001110";
Trees_din <= "00000100000000000011000100000100";
wait for Clk_period;
Addr <= "1001010001111";
Trees_din <= "00000000001011010100101001100001";
wait for Clk_period;
Addr <= "1001010010000";
Trees_din <= "00000000000110110100101001100001";
wait for Clk_period;
Addr <= "1001010010001";
Trees_din <= "00000100000000000010100000001000";
wait for Clk_period;
Addr <= "1001010010010";
Trees_din <= "00000010000000000011001100000100";
wait for Clk_period;
Addr <= "1001010010011";
Trees_din <= "00000000010001010100101001100001";
wait for Clk_period;
Addr <= "1001010010100";
Trees_din <= "00000000001110010100101001100001";
wait for Clk_period;
Addr <= "1001010010101";
Trees_din <= "00000001000000000001001100000100";
wait for Clk_period;
Addr <= "1001010010110";
Trees_din <= "00000000010110110100101001100001";
wait for Clk_period;
Addr <= "1001010010111";
Trees_din <= "00000000010110010100101001100001";
wait for Clk_period;



----------tree 37-------------------

Addr <= "1001010011000";
Trees_din <= "00000010000000000010111110000000";
wait for Clk_period;
Addr <= "1001010011001";
Trees_din <= "00000001000000000100000101000000";
wait for Clk_period;
Addr <= "1001010011010";
Trees_din <= "00000000000000000010000000100000";
wait for Clk_period;
Addr <= "1001010011011";
Trees_din <= "00000001000000000100111100010000";
wait for Clk_period;
Addr <= "1001010011100";
Trees_din <= "00000010000000000001000100001000";
wait for Clk_period;
Addr <= "1001010011101";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "1001010011110";
Trees_din <= "00000000010100110100110001011101";
wait for Clk_period;
Addr <= "1001010011111";
Trees_din <= "00000000000011100100110001011101";
wait for Clk_period;
Addr <= "1001010100000";
Trees_din <= "00000010000000000010000000000100";
wait for Clk_period;
Addr <= "1001010100001";
Trees_din <= "00000000001100010100110001011101";
wait for Clk_period;
Addr <= "1001010100010";
Trees_din <= "00000000000101100100110001011101";
wait for Clk_period;
Addr <= "1001010100011";
Trees_din <= "00000111000000000010011000001000";
wait for Clk_period;
Addr <= "1001010100100";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "1001010100101";
Trees_din <= "00000000010011110100110001011101";
wait for Clk_period;
Addr <= "1001010100110";
Trees_din <= "00000000010010100100110001011101";
wait for Clk_period;
Addr <= "1001010100111";
Trees_din <= "00000011000000000101010100000100";
wait for Clk_period;
Addr <= "1001010101000";
Trees_din <= "00000000000111110100110001011101";
wait for Clk_period;
Addr <= "1001010101001";
Trees_din <= "00000000010011100100110001011101";
wait for Clk_period;
Addr <= "1001010101010";
Trees_din <= "00000001000000000011100000010000";
wait for Clk_period;
Addr <= "1001010101011";
Trees_din <= "00000001000000000000111100001000";
wait for Clk_period;
Addr <= "1001010101100";
Trees_din <= "00000000000000000011100000000100";
wait for Clk_period;
Addr <= "1001010101101";
Trees_din <= "00000000001010110100110001011101";
wait for Clk_period;
Addr <= "1001010101110";
Trees_din <= "00000000010110100100110001011101";
wait for Clk_period;
Addr <= "1001010101111";
Trees_din <= "00000110000000000101110100000100";
wait for Clk_period;
Addr <= "1001010110000";
Trees_din <= "00000000010010100100110001011101";
wait for Clk_period;
Addr <= "1001010110001";
Trees_din <= "00000000001010110100110001011101";
wait for Clk_period;
Addr <= "1001010110010";
Trees_din <= "00000001000000000001110000001000";
wait for Clk_period;
Addr <= "1001010110011";
Trees_din <= "00000001000000000010111000000100";
wait for Clk_period;
Addr <= "1001010110100";
Trees_din <= "00000000010101010100110001011101";
wait for Clk_period;
Addr <= "1001010110101";
Trees_din <= "00000000000110100100110001011101";
wait for Clk_period;
Addr <= "1001010110110";
Trees_din <= "00000000000000000011000000000100";
wait for Clk_period;
Addr <= "1001010110111";
Trees_din <= "00000000010111100100110001011101";
wait for Clk_period;
Addr <= "1001010111000";
Trees_din <= "00000000001001010100110001011101";
wait for Clk_period;
Addr <= "1001010111001";
Trees_din <= "00000010000000000011100000100000";
wait for Clk_period;
Addr <= "1001010111010";
Trees_din <= "00000111000000000011001100010000";
wait for Clk_period;
Addr <= "1001010111011";
Trees_din <= "00000001000000000101110100001000";
wait for Clk_period;
Addr <= "1001010111100";
Trees_din <= "00000111000000000000111000000100";
wait for Clk_period;
Addr <= "1001010111101";
Trees_din <= "00000000011000010100110001011101";
wait for Clk_period;
Addr <= "1001010111110";
Trees_din <= "00000000000000010100110001011101";
wait for Clk_period;
Addr <= "1001010111111";
Trees_din <= "00000111000000000011111000000100";
wait for Clk_period;
Addr <= "1001011000000";
Trees_din <= "00000000000011000100110001011101";
wait for Clk_period;
Addr <= "1001011000001";
Trees_din <= "00000000000000100100110001011101";
wait for Clk_period;
Addr <= "1001011000010";
Trees_din <= "00000010000000000100011100001000";
wait for Clk_period;
Addr <= "1001011000011";
Trees_din <= "00000110000000000010011100000100";
wait for Clk_period;
Addr <= "1001011000100";
Trees_din <= "00000000001100100100110001011101";
wait for Clk_period;
Addr <= "1001011000101";
Trees_din <= "00000000001100000100110001011101";
wait for Clk_period;
Addr <= "1001011000110";
Trees_din <= "00000011000000000001001100000100";
wait for Clk_period;
Addr <= "1001011000111";
Trees_din <= "00000000001010110100110001011101";
wait for Clk_period;
Addr <= "1001011001000";
Trees_din <= "00000000001000100100110001011101";
wait for Clk_period;
Addr <= "1001011001001";
Trees_din <= "00000110000000000010101000010000";
wait for Clk_period;
Addr <= "1001011001010";
Trees_din <= "00000011000000000001110100001000";
wait for Clk_period;
Addr <= "1001011001011";
Trees_din <= "00000100000000000100110100000100";
wait for Clk_period;
Addr <= "1001011001100";
Trees_din <= "00000000010010000100110001011101";
wait for Clk_period;
Addr <= "1001011001101";
Trees_din <= "00000000010101110100110001011101";
wait for Clk_period;
Addr <= "1001011001110";
Trees_din <= "00000001000000000000010000000100";
wait for Clk_period;
Addr <= "1001011001111";
Trees_din <= "00000000001111100100110001011101";
wait for Clk_period;
Addr <= "1001011010000";
Trees_din <= "00000000010001000100110001011101";
wait for Clk_period;
Addr <= "1001011010001";
Trees_din <= "00000101000000000100011000001000";
wait for Clk_period;
Addr <= "1001011010010";
Trees_din <= "00000010000000000001111100000100";
wait for Clk_period;
Addr <= "1001011010011";
Trees_din <= "00000000010001100100110001011101";
wait for Clk_period;
Addr <= "1001011010100";
Trees_din <= "00000000001000000100110001011101";
wait for Clk_period;
Addr <= "1001011010101";
Trees_din <= "00000111000000000001100100000100";
wait for Clk_period;
Addr <= "1001011010110";
Trees_din <= "00000000011000000100110001011101";
wait for Clk_period;
Addr <= "1001011010111";
Trees_din <= "00000000010100110100110001011101";
wait for Clk_period;
Addr <= "1001011011000";
Trees_din <= "00000110000000000000111001000000";
wait for Clk_period;
Addr <= "1001011011001";
Trees_din <= "00000101000000000010110100100000";
wait for Clk_period;
Addr <= "1001011011010";
Trees_din <= "00000100000000000010011100010000";
wait for Clk_period;
Addr <= "1001011011011";
Trees_din <= "00000111000000000001111100001000";
wait for Clk_period;
Addr <= "1001011011100";
Trees_din <= "00000011000000000010100100000100";
wait for Clk_period;
Addr <= "1001011011101";
Trees_din <= "00000000000001100100110001011101";
wait for Clk_period;
Addr <= "1001011011110";
Trees_din <= "00000000000111100100110001011101";
wait for Clk_period;
Addr <= "1001011011111";
Trees_din <= "00000100000000000011100100000100";
wait for Clk_period;
Addr <= "1001011100000";
Trees_din <= "00000000001000110100110001011101";
wait for Clk_period;
Addr <= "1001011100001";
Trees_din <= "00000000010100000100110001011101";
wait for Clk_period;
Addr <= "1001011100010";
Trees_din <= "00000010000000000110000000001000";
wait for Clk_period;
Addr <= "1001011100011";
Trees_din <= "00000111000000000101010100000100";
wait for Clk_period;
Addr <= "1001011100100";
Trees_din <= "00000000000110100100110001011101";
wait for Clk_period;
Addr <= "1001011100101";
Trees_din <= "00000000001010010100110001011101";
wait for Clk_period;
Addr <= "1001011100110";
Trees_din <= "00000110000000000011001100000100";
wait for Clk_period;
Addr <= "1001011100111";
Trees_din <= "00000000010111000100110001011101";
wait for Clk_period;
Addr <= "1001011101000";
Trees_din <= "00000000000011100100110001011101";
wait for Clk_period;
Addr <= "1001011101001";
Trees_din <= "00000001000000000011101100010000";
wait for Clk_period;
Addr <= "1001011101010";
Trees_din <= "00000111000000000011101000001000";
wait for Clk_period;
Addr <= "1001011101011";
Trees_din <= "00000000000000000000010100000100";
wait for Clk_period;
Addr <= "1001011101100";
Trees_din <= "00000000000100010100110001011101";
wait for Clk_period;
Addr <= "1001011101101";
Trees_din <= "00000000010010110100110001011101";
wait for Clk_period;
Addr <= "1001011101110";
Trees_din <= "00000000000000000011001100000100";
wait for Clk_period;
Addr <= "1001011101111";
Trees_din <= "00000000000000110100110001011101";
wait for Clk_period;
Addr <= "1001011110000";
Trees_din <= "00000000010100000100110001011101";
wait for Clk_period;
Addr <= "1001011110001";
Trees_din <= "00000101000000000011001000001000";
wait for Clk_period;
Addr <= "1001011110010";
Trees_din <= "00000101000000000011110100000100";
wait for Clk_period;
Addr <= "1001011110011";
Trees_din <= "00000000010011010100110001011101";
wait for Clk_period;
Addr <= "1001011110100";
Trees_din <= "00000000010110000100110001011101";
wait for Clk_period;
Addr <= "1001011110101";
Trees_din <= "00000011000000000101011100000100";
wait for Clk_period;
Addr <= "1001011110110";
Trees_din <= "00000000000101110100110001011101";
wait for Clk_period;
Addr <= "1001011110111";
Trees_din <= "00000000010100010100110001011101";
wait for Clk_period;
Addr <= "1001011111000";
Trees_din <= "00000011000000000001000100100000";
wait for Clk_period;
Addr <= "1001011111001";
Trees_din <= "00000100000000000011111100010000";
wait for Clk_period;
Addr <= "1001011111010";
Trees_din <= "00000100000000000000000100001000";
wait for Clk_period;
Addr <= "1001011111011";
Trees_din <= "00000000000000000101001100000100";
wait for Clk_period;
Addr <= "1001011111100";
Trees_din <= "00000000001011000100110001011101";
wait for Clk_period;
Addr <= "1001011111101";
Trees_din <= "00000000000000010100110001011101";
wait for Clk_period;
Addr <= "1001011111110";
Trees_din <= "00000000000000000010111000000100";
wait for Clk_period;
Addr <= "1001011111111";
Trees_din <= "00000000010111100100110001011101";
wait for Clk_period;
Addr <= "1001100000000";
Trees_din <= "00000000000101110100110001011101";
wait for Clk_period;
Addr <= "1001100000001";
Trees_din <= "00000100000000000010000000001000";
wait for Clk_period;
Addr <= "1001100000010";
Trees_din <= "00000110000000000010110100000100";
wait for Clk_period;
Addr <= "1001100000011";
Trees_din <= "00000000010100000100110001011101";
wait for Clk_period;
Addr <= "1001100000100";
Trees_din <= "00000000010110100100110001011101";
wait for Clk_period;
Addr <= "1001100000101";
Trees_din <= "00000001000000000001100100000100";
wait for Clk_period;
Addr <= "1001100000110";
Trees_din <= "00000000010000010100110001011101";
wait for Clk_period;
Addr <= "1001100000111";
Trees_din <= "00000000010011110100110001011101";
wait for Clk_period;
Addr <= "1001100001000";
Trees_din <= "00000001000000000000000000010000";
wait for Clk_period;
Addr <= "1001100001001";
Trees_din <= "00000000000000000000010000001000";
wait for Clk_period;
Addr <= "1001100001010";
Trees_din <= "00000010000000000000010000000100";
wait for Clk_period;
Addr <= "1001100001011";
Trees_din <= "00000000010010110100110001011101";
wait for Clk_period;
Addr <= "1001100001100";
Trees_din <= "00000000000000110100110001011101";
wait for Clk_period;
Addr <= "1001100001101";
Trees_din <= "00000011000000000010001000000100";
wait for Clk_period;
Addr <= "1001100001110";
Trees_din <= "00000000001100000100110001011101";
wait for Clk_period;
Addr <= "1001100001111";
Trees_din <= "00000000010101110100110001011101";
wait for Clk_period;
Addr <= "1001100010000";
Trees_din <= "00000101000000000101010000001000";
wait for Clk_period;
Addr <= "1001100010001";
Trees_din <= "00000000000000000001000100000100";
wait for Clk_period;
Addr <= "1001100010010";
Trees_din <= "00000000010101110100110001011101";
wait for Clk_period;
Addr <= "1001100010011";
Trees_din <= "00000000000101110100110001011101";
wait for Clk_period;
Addr <= "1001100010100";
Trees_din <= "00000011000000000100111000000100";
wait for Clk_period;
Addr <= "1001100010101";
Trees_din <= "00000000000101100100110001011101";
wait for Clk_period;
Addr <= "1001100010110";
Trees_din <= "00000000011000000100110001011101";
wait for Clk_period;



----------tree 38-------------------

Addr <= "1001100010111";
Trees_din <= "00000000000000000001011010000000";
wait for Clk_period;
Addr <= "1001100011000";
Trees_din <= "00000000000000000011000001000000";
wait for Clk_period;
Addr <= "1001100011001";
Trees_din <= "00000001000000000000010000100000";
wait for Clk_period;
Addr <= "1001100011010";
Trees_din <= "00000101000000000011110100010000";
wait for Clk_period;
Addr <= "1001100011011";
Trees_din <= "00000000000000000101110100001000";
wait for Clk_period;
Addr <= "1001100011100";
Trees_din <= "00000100000000000100010100000100";
wait for Clk_period;
Addr <= "1001100011101";
Trees_din <= "00000000001111100100111001011001";
wait for Clk_period;
Addr <= "1001100011110";
Trees_din <= "00000000011001000100111001011001";
wait for Clk_period;
Addr <= "1001100011111";
Trees_din <= "00000101000000000011011000000100";
wait for Clk_period;
Addr <= "1001100100000";
Trees_din <= "00000000000111010100111001011001";
wait for Clk_period;
Addr <= "1001100100001";
Trees_din <= "00000000001000100100111001011001";
wait for Clk_period;
Addr <= "1001100100010";
Trees_din <= "00000001000000000001101100001000";
wait for Clk_period;
Addr <= "1001100100011";
Trees_din <= "00000011000000000101101100000100";
wait for Clk_period;
Addr <= "1001100100100";
Trees_din <= "00000000011000100100111001011001";
wait for Clk_period;
Addr <= "1001100100101";
Trees_din <= "00000000000110000100111001011001";
wait for Clk_period;
Addr <= "1001100100110";
Trees_din <= "00000101000000000101110100000100";
wait for Clk_period;
Addr <= "1001100100111";
Trees_din <= "00000000000111010100111001011001";
wait for Clk_period;
Addr <= "1001100101000";
Trees_din <= "00000000001101000100111001011001";
wait for Clk_period;
Addr <= "1001100101001";
Trees_din <= "00000101000000000100011000010000";
wait for Clk_period;
Addr <= "1001100101010";
Trees_din <= "00000000000000000000111100001000";
wait for Clk_period;
Addr <= "1001100101011";
Trees_din <= "00000000000000000001100100000100";
wait for Clk_period;
Addr <= "1001100101100";
Trees_din <= "00000000001110000100111001011001";
wait for Clk_period;
Addr <= "1001100101101";
Trees_din <= "00000000001011110100111001011001";
wait for Clk_period;
Addr <= "1001100101110";
Trees_din <= "00000010000000000001100000000100";
wait for Clk_period;
Addr <= "1001100101111";
Trees_din <= "00000000000110100100111001011001";
wait for Clk_period;
Addr <= "1001100110000";
Trees_din <= "00000000001101000100111001011001";
wait for Clk_period;
Addr <= "1001100110001";
Trees_din <= "00000011000000000001111000001000";
wait for Clk_period;
Addr <= "1001100110010";
Trees_din <= "00000010000000000000110000000100";
wait for Clk_period;
Addr <= "1001100110011";
Trees_din <= "00000000010001000100111001011001";
wait for Clk_period;
Addr <= "1001100110100";
Trees_din <= "00000000001110010100111001011001";
wait for Clk_period;
Addr <= "1001100110101";
Trees_din <= "00000011000000000010100000000100";
wait for Clk_period;
Addr <= "1001100110110";
Trees_din <= "00000000000110100100111001011001";
wait for Clk_period;
Addr <= "1001100110111";
Trees_din <= "00000000001101010100111001011001";
wait for Clk_period;
Addr <= "1001100111000";
Trees_din <= "00000010000000000001010100100000";
wait for Clk_period;
Addr <= "1001100111001";
Trees_din <= "00000101000000000100010000010000";
wait for Clk_period;
Addr <= "1001100111010";
Trees_din <= "00000100000000000010010000001000";
wait for Clk_period;
Addr <= "1001100111011";
Trees_din <= "00000110000000000000100000000100";
wait for Clk_period;
Addr <= "1001100111100";
Trees_din <= "00000000001111000100111001011001";
wait for Clk_period;
Addr <= "1001100111101";
Trees_din <= "00000000001000100100111001011001";
wait for Clk_period;
Addr <= "1001100111110";
Trees_din <= "00000110000000000100111000000100";
wait for Clk_period;
Addr <= "1001100111111";
Trees_din <= "00000000000001100100111001011001";
wait for Clk_period;
Addr <= "1001101000000";
Trees_din <= "00000000000000000100111001011001";
wait for Clk_period;
Addr <= "1001101000001";
Trees_din <= "00000001000000000101110000001000";
wait for Clk_period;
Addr <= "1001101000010";
Trees_din <= "00000011000000000011100000000100";
wait for Clk_period;
Addr <= "1001101000011";
Trees_din <= "00000000001011110100111001011001";
wait for Clk_period;
Addr <= "1001101000100";
Trees_din <= "00000000010011100100111001011001";
wait for Clk_period;
Addr <= "1001101000101";
Trees_din <= "00000110000000000100010100000100";
wait for Clk_period;
Addr <= "1001101000110";
Trees_din <= "00000000010101010100111001011001";
wait for Clk_period;
Addr <= "1001101000111";
Trees_din <= "00000000010110000100111001011001";
wait for Clk_period;
Addr <= "1001101001000";
Trees_din <= "00000001000000000011000100010000";
wait for Clk_period;
Addr <= "1001101001001";
Trees_din <= "00000110000000000001011100001000";
wait for Clk_period;
Addr <= "1001101001010";
Trees_din <= "00000111000000000001100000000100";
wait for Clk_period;
Addr <= "1001101001011";
Trees_din <= "00000000010000010100111001011001";
wait for Clk_period;
Addr <= "1001101001100";
Trees_din <= "00000000001010000100111001011001";
wait for Clk_period;
Addr <= "1001101001101";
Trees_din <= "00000011000000000000011100000100";
wait for Clk_period;
Addr <= "1001101001110";
Trees_din <= "00000000010101110100111001011001";
wait for Clk_period;
Addr <= "1001101001111";
Trees_din <= "00000000001110100100111001011001";
wait for Clk_period;
Addr <= "1001101010000";
Trees_din <= "00000111000000000000110000001000";
wait for Clk_period;
Addr <= "1001101010001";
Trees_din <= "00000011000000000100001000000100";
wait for Clk_period;
Addr <= "1001101010010";
Trees_din <= "00000000001100110100111001011001";
wait for Clk_period;
Addr <= "1001101010011";
Trees_din <= "00000000000111000100111001011001";
wait for Clk_period;
Addr <= "1001101010100";
Trees_din <= "00000110000000000101111000000100";
wait for Clk_period;
Addr <= "1001101010101";
Trees_din <= "00000000001110100100111001011001";
wait for Clk_period;
Addr <= "1001101010110";
Trees_din <= "00000000010101110100111001011001";
wait for Clk_period;
Addr <= "1001101010111";
Trees_din <= "00000000000000000101111001000000";
wait for Clk_period;
Addr <= "1001101011000";
Trees_din <= "00000001000000000100011000100000";
wait for Clk_period;
Addr <= "1001101011001";
Trees_din <= "00000110000000000000011000010000";
wait for Clk_period;
Addr <= "1001101011010";
Trees_din <= "00000001000000000001000000001000";
wait for Clk_period;
Addr <= "1001101011011";
Trees_din <= "00000001000000000011011100000100";
wait for Clk_period;
Addr <= "1001101011100";
Trees_din <= "00000000010100000100111001011001";
wait for Clk_period;
Addr <= "1001101011101";
Trees_din <= "00000000000000010100111001011001";
wait for Clk_period;
Addr <= "1001101011110";
Trees_din <= "00000110000000000000101000000100";
wait for Clk_period;
Addr <= "1001101011111";
Trees_din <= "00000000000101010100111001011001";
wait for Clk_period;
Addr <= "1001101100000";
Trees_din <= "00000000010110100100111001011001";
wait for Clk_period;
Addr <= "1001101100001";
Trees_din <= "00000110000000000000110100001000";
wait for Clk_period;
Addr <= "1001101100010";
Trees_din <= "00000101000000000010010100000100";
wait for Clk_period;
Addr <= "1001101100011";
Trees_din <= "00000000000011000100111001011001";
wait for Clk_period;
Addr <= "1001101100100";
Trees_din <= "00000000000011000100111001011001";
wait for Clk_period;
Addr <= "1001101100101";
Trees_din <= "00000001000000000001110000000100";
wait for Clk_period;
Addr <= "1001101100110";
Trees_din <= "00000000000010110100111001011001";
wait for Clk_period;
Addr <= "1001101100111";
Trees_din <= "00000000001100100100111001011001";
wait for Clk_period;
Addr <= "1001101101000";
Trees_din <= "00000010000000000000011100010000";
wait for Clk_period;
Addr <= "1001101101001";
Trees_din <= "00000000000000000101101000001000";
wait for Clk_period;
Addr <= "1001101101010";
Trees_din <= "00000100000000000011110000000100";
wait for Clk_period;
Addr <= "1001101101011";
Trees_din <= "00000000001111000100111001011001";
wait for Clk_period;
Addr <= "1001101101100";
Trees_din <= "00000000001001000100111001011001";
wait for Clk_period;
Addr <= "1001101101101";
Trees_din <= "00000011000000000010101000000100";
wait for Clk_period;
Addr <= "1001101101110";
Trees_din <= "00000000000001010100111001011001";
wait for Clk_period;
Addr <= "1001101101111";
Trees_din <= "00000000000010100100111001011001";
wait for Clk_period;
Addr <= "1001101110000";
Trees_din <= "00000101000000000000110000001000";
wait for Clk_period;
Addr <= "1001101110001";
Trees_din <= "00000011000000000001111100000100";
wait for Clk_period;
Addr <= "1001101110010";
Trees_din <= "00000000011000000100111001011001";
wait for Clk_period;
Addr <= "1001101110011";
Trees_din <= "00000000001011110100111001011001";
wait for Clk_period;
Addr <= "1001101110100";
Trees_din <= "00000010000000000000011100000100";
wait for Clk_period;
Addr <= "1001101110101";
Trees_din <= "00000000010001100100111001011001";
wait for Clk_period;
Addr <= "1001101110110";
Trees_din <= "00000000010010010100111001011001";
wait for Clk_period;
Addr <= "1001101110111";
Trees_din <= "00000010000000000101010000100000";
wait for Clk_period;
Addr <= "1001101111000";
Trees_din <= "00000010000000000001110100010000";
wait for Clk_period;
Addr <= "1001101111001";
Trees_din <= "00000000000000000000110100001000";
wait for Clk_period;
Addr <= "1001101111010";
Trees_din <= "00000000000000000010111000000100";
wait for Clk_period;
Addr <= "1001101111011";
Trees_din <= "00000000010110100100111001011001";
wait for Clk_period;
Addr <= "1001101111100";
Trees_din <= "00000000000100100100111001011001";
wait for Clk_period;
Addr <= "1001101111101";
Trees_din <= "00000010000000000001001000000100";
wait for Clk_period;
Addr <= "1001101111110";
Trees_din <= "00000000001010000100111001011001";
wait for Clk_period;
Addr <= "1001101111111";
Trees_din <= "00000000010111110100111001011001";
wait for Clk_period;
Addr <= "1001110000000";
Trees_din <= "00000111000000000010101100001000";
wait for Clk_period;
Addr <= "1001110000001";
Trees_din <= "00000000000000000101001100000100";
wait for Clk_period;
Addr <= "1001110000010";
Trees_din <= "00000000001010100100111001011001";
wait for Clk_period;
Addr <= "1001110000011";
Trees_din <= "00000000011001000100111001011001";
wait for Clk_period;
Addr <= "1001110000100";
Trees_din <= "00000111000000000000100100000100";
wait for Clk_period;
Addr <= "1001110000101";
Trees_din <= "00000000010111100100111001011001";
wait for Clk_period;
Addr <= "1001110000110";
Trees_din <= "00000000000101110100111001011001";
wait for Clk_period;
Addr <= "1001110000111";
Trees_din <= "00000101000000000101001000010000";
wait for Clk_period;
Addr <= "1001110001000";
Trees_din <= "00000010000000000000000000001000";
wait for Clk_period;
Addr <= "1001110001001";
Trees_din <= "00000011000000000010111000000100";
wait for Clk_period;
Addr <= "1001110001010";
Trees_din <= "00000000010100100100111001011001";
wait for Clk_period;
Addr <= "1001110001011";
Trees_din <= "00000000011000000100111001011001";
wait for Clk_period;
Addr <= "1001110001100";
Trees_din <= "00000001000000000000111000000100";
wait for Clk_period;
Addr <= "1001110001101";
Trees_din <= "00000000010011010100111001011001";
wait for Clk_period;
Addr <= "1001110001110";
Trees_din <= "00000000000000000100111001011001";
wait for Clk_period;
Addr <= "1001110001111";
Trees_din <= "00000010000000000001110100001000";
wait for Clk_period;
Addr <= "1001110010000";
Trees_din <= "00000011000000000010001000000100";
wait for Clk_period;
Addr <= "1001110010001";
Trees_din <= "00000000001111000100111001011001";
wait for Clk_period;
Addr <= "1001110010010";
Trees_din <= "00000000010010000100111001011001";
wait for Clk_period;
Addr <= "1001110010011";
Trees_din <= "00000001000000000000110100000100";
wait for Clk_period;
Addr <= "1001110010100";
Trees_din <= "00000000010111000100111001011001";
wait for Clk_period;
Addr <= "1001110010101";
Trees_din <= "00000000010111010100111001011001";
wait for Clk_period;



----------tree 39-------------------

Addr <= "1001110010110";
Trees_din <= "00000001000000000100011010000000";
wait for Clk_period;
Addr <= "1001110010111";
Trees_din <= "00000101000000000100111101000000";
wait for Clk_period;
Addr <= "1001110011000";
Trees_din <= "00000110000000000000101100100000";
wait for Clk_period;
Addr <= "1001110011001";
Trees_din <= "00000101000000000000011000010000";
wait for Clk_period;
Addr <= "1001110011010";
Trees_din <= "00000110000000000001011000001000";
wait for Clk_period;
Addr <= "1001110011011";
Trees_din <= "00000011000000000101110000000100";
wait for Clk_period;
Addr <= "1001110011100";
Trees_din <= "00000000010001110101000001010101";
wait for Clk_period;
Addr <= "1001110011101";
Trees_din <= "00000000010100110101000001010101";
wait for Clk_period;
Addr <= "1001110011110";
Trees_din <= "00000001000000000001111000000100";
wait for Clk_period;
Addr <= "1001110011111";
Trees_din <= "00000000001101100101000001010101";
wait for Clk_period;
Addr <= "1001110100000";
Trees_din <= "00000000000101100101000001010101";
wait for Clk_period;
Addr <= "1001110100001";
Trees_din <= "00000101000000000001111000001000";
wait for Clk_period;
Addr <= "1001110100010";
Trees_din <= "00000101000000000100010100000100";
wait for Clk_period;
Addr <= "1001110100011";
Trees_din <= "00000000010101100101000001010101";
wait for Clk_period;
Addr <= "1001110100100";
Trees_din <= "00000000001111100101000001010101";
wait for Clk_period;
Addr <= "1001110100101";
Trees_din <= "00000011000000000010111000000100";
wait for Clk_period;
Addr <= "1001110100110";
Trees_din <= "00000000010100010101000001010101";
wait for Clk_period;
Addr <= "1001110100111";
Trees_din <= "00000000001011110101000001010101";
wait for Clk_period;
Addr <= "1001110101000";
Trees_din <= "00000000000000000000000100010000";
wait for Clk_period;
Addr <= "1001110101001";
Trees_din <= "00000111000000000010010100001000";
wait for Clk_period;
Addr <= "1001110101010";
Trees_din <= "00000011000000000101011100000100";
wait for Clk_period;
Addr <= "1001110101011";
Trees_din <= "00000000010100100101000001010101";
wait for Clk_period;
Addr <= "1001110101100";
Trees_din <= "00000000010010010101000001010101";
wait for Clk_period;
Addr <= "1001110101101";
Trees_din <= "00000101000000000011000000000100";
wait for Clk_period;
Addr <= "1001110101110";
Trees_din <= "00000000000111000101000001010101";
wait for Clk_period;
Addr <= "1001110101111";
Trees_din <= "00000000001100000101000001010101";
wait for Clk_period;
Addr <= "1001110110000";
Trees_din <= "00000000000000000000010100001000";
wait for Clk_period;
Addr <= "1001110110001";
Trees_din <= "00000100000000000100011000000100";
wait for Clk_period;
Addr <= "1001110110010";
Trees_din <= "00000000000100100101000001010101";
wait for Clk_period;
Addr <= "1001110110011";
Trees_din <= "00000000001000000101000001010101";
wait for Clk_period;
Addr <= "1001110110100";
Trees_din <= "00000100000000000001110000000100";
wait for Clk_period;
Addr <= "1001110110101";
Trees_din <= "00000000000011100101000001010101";
wait for Clk_period;
Addr <= "1001110110110";
Trees_din <= "00000000001010110101000001010101";
wait for Clk_period;
Addr <= "1001110110111";
Trees_din <= "00000110000000000000100100100000";
wait for Clk_period;
Addr <= "1001110111000";
Trees_din <= "00000000000000000010010100010000";
wait for Clk_period;
Addr <= "1001110111001";
Trees_din <= "00000000000000000101010000001000";
wait for Clk_period;
Addr <= "1001110111010";
Trees_din <= "00000011000000000011101000000100";
wait for Clk_period;
Addr <= "1001110111011";
Trees_din <= "00000000001010000101000001010101";
wait for Clk_period;
Addr <= "1001110111100";
Trees_din <= "00000000010010010101000001010101";
wait for Clk_period;
Addr <= "1001110111101";
Trees_din <= "00000101000000000100000000000100";
wait for Clk_period;
Addr <= "1001110111110";
Trees_din <= "00000000010111010101000001010101";
wait for Clk_period;
Addr <= "1001110111111";
Trees_din <= "00000000001101110101000001010101";
wait for Clk_period;
Addr <= "1001111000000";
Trees_din <= "00000010000000000001100100001000";
wait for Clk_period;
Addr <= "1001111000001";
Trees_din <= "00000101000000000000001000000100";
wait for Clk_period;
Addr <= "1001111000010";
Trees_din <= "00000000001110000101000001010101";
wait for Clk_period;
Addr <= "1001111000011";
Trees_din <= "00000000010001110101000001010101";
wait for Clk_period;
Addr <= "1001111000100";
Trees_din <= "00000001000000000100000000000100";
wait for Clk_period;
Addr <= "1001111000101";
Trees_din <= "00000000000011100101000001010101";
wait for Clk_period;
Addr <= "1001111000110";
Trees_din <= "00000000010010010101000001010101";
wait for Clk_period;
Addr <= "1001111000111";
Trees_din <= "00000001000000000011001100010000";
wait for Clk_period;
Addr <= "1001111001000";
Trees_din <= "00000111000000000011011000001000";
wait for Clk_period;
Addr <= "1001111001001";
Trees_din <= "00000000000000000101010100000100";
wait for Clk_period;
Addr <= "1001111001010";
Trees_din <= "00000000010001000101000001010101";
wait for Clk_period;
Addr <= "1001111001011";
Trees_din <= "00000000001100000101000001010101";
wait for Clk_period;
Addr <= "1001111001100";
Trees_din <= "00000101000000000101010100000100";
wait for Clk_period;
Addr <= "1001111001101";
Trees_din <= "00000000010001010101000001010101";
wait for Clk_period;
Addr <= "1001111001110";
Trees_din <= "00000000010000010101000001010101";
wait for Clk_period;
Addr <= "1001111001111";
Trees_din <= "00000110000000000001001100001000";
wait for Clk_period;
Addr <= "1001111010000";
Trees_din <= "00000000000000000101110000000100";
wait for Clk_period;
Addr <= "1001111010001";
Trees_din <= "00000000001011010101000001010101";
wait for Clk_period;
Addr <= "1001111010010";
Trees_din <= "00000000001010000101000001010101";
wait for Clk_period;
Addr <= "1001111010011";
Trees_din <= "00000001000000000001000000000100";
wait for Clk_period;
Addr <= "1001111010100";
Trees_din <= "00000000010011010101000001010101";
wait for Clk_period;
Addr <= "1001111010101";
Trees_din <= "00000000000110010101000001010101";
wait for Clk_period;
Addr <= "1001111010110";
Trees_din <= "00000100000000000001011001000000";
wait for Clk_period;
Addr <= "1001111010111";
Trees_din <= "00000100000000000100000000100000";
wait for Clk_period;
Addr <= "1001111011000";
Trees_din <= "00000011000000000010110100010000";
wait for Clk_period;
Addr <= "1001111011001";
Trees_din <= "00000010000000000000010100001000";
wait for Clk_period;
Addr <= "1001111011010";
Trees_din <= "00000011000000000100111100000100";
wait for Clk_period;
Addr <= "1001111011011";
Trees_din <= "00000000001000110101000001010101";
wait for Clk_period;
Addr <= "1001111011100";
Trees_din <= "00000000010000010101000001010101";
wait for Clk_period;
Addr <= "1001111011101";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "1001111011110";
Trees_din <= "00000000000101010101000001010101";
wait for Clk_period;
Addr <= "1001111011111";
Trees_din <= "00000000001111100101000001010101";
wait for Clk_period;
Addr <= "1001111100000";
Trees_din <= "00000001000000000010101100001000";
wait for Clk_period;
Addr <= "1001111100001";
Trees_din <= "00000001000000000011000000000100";
wait for Clk_period;
Addr <= "1001111100010";
Trees_din <= "00000000010010100101000001010101";
wait for Clk_period;
Addr <= "1001111100011";
Trees_din <= "00000000011000100101000001010101";
wait for Clk_period;
Addr <= "1001111100100";
Trees_din <= "00000001000000000010110000000100";
wait for Clk_period;
Addr <= "1001111100101";
Trees_din <= "00000000010011100101000001010101";
wait for Clk_period;
Addr <= "1001111100110";
Trees_din <= "00000000000011010101000001010101";
wait for Clk_period;
Addr <= "1001111100111";
Trees_din <= "00000110000000000101001100010000";
wait for Clk_period;
Addr <= "1001111101000";
Trees_din <= "00000001000000000001011000001000";
wait for Clk_period;
Addr <= "1001111101001";
Trees_din <= "00000101000000000000010100000100";
wait for Clk_period;
Addr <= "1001111101010";
Trees_din <= "00000000001000110101000001010101";
wait for Clk_period;
Addr <= "1001111101011";
Trees_din <= "00000000001101000101000001010101";
wait for Clk_period;
Addr <= "1001111101100";
Trees_din <= "00000100000000000100010000000100";
wait for Clk_period;
Addr <= "1001111101101";
Trees_din <= "00000000010000000101000001010101";
wait for Clk_period;
Addr <= "1001111101110";
Trees_din <= "00000000000010010101000001010101";
wait for Clk_period;
Addr <= "1001111101111";
Trees_din <= "00000000000000000101100100001000";
wait for Clk_period;
Addr <= "1001111110000";
Trees_din <= "00000011000000000011110100000100";
wait for Clk_period;
Addr <= "1001111110001";
Trees_din <= "00000000010110010101000001010101";
wait for Clk_period;
Addr <= "1001111110010";
Trees_din <= "00000000001001000101000001010101";
wait for Clk_period;
Addr <= "1001111110011";
Trees_din <= "00000100000000000000000000000100";
wait for Clk_period;
Addr <= "1001111110100";
Trees_din <= "00000000010111000101000001010101";
wait for Clk_period;
Addr <= "1001111110101";
Trees_din <= "00000000001000100101000001010101";
wait for Clk_period;
Addr <= "1001111110110";
Trees_din <= "00000110000000000011010100100000";
wait for Clk_period;
Addr <= "1001111110111";
Trees_din <= "00000001000000000001011000010000";
wait for Clk_period;
Addr <= "1001111111000";
Trees_din <= "00000000000000000001010100001000";
wait for Clk_period;
Addr <= "1001111111001";
Trees_din <= "00000110000000000000101000000100";
wait for Clk_period;
Addr <= "1001111111010";
Trees_din <= "00000000010110010101000001010101";
wait for Clk_period;
Addr <= "1001111111011";
Trees_din <= "00000000001010110101000001010101";
wait for Clk_period;
Addr <= "1001111111100";
Trees_din <= "00000001000000000011111000000100";
wait for Clk_period;
Addr <= "1001111111101";
Trees_din <= "00000000001101000101000001010101";
wait for Clk_period;
Addr <= "1001111111110";
Trees_din <= "00000000010101110101000001010101";
wait for Clk_period;
Addr <= "1001111111111";
Trees_din <= "00000100000000000011100000001000";
wait for Clk_period;
Addr <= "1010000000000";
Trees_din <= "00000111000000000011101000000100";
wait for Clk_period;
Addr <= "1010000000001";
Trees_din <= "00000000000011110101000001010101";
wait for Clk_period;
Addr <= "1010000000010";
Trees_din <= "00000000001011000101000001010101";
wait for Clk_period;
Addr <= "1010000000011";
Trees_din <= "00000001000000000100101000000100";
wait for Clk_period;
Addr <= "1010000000100";
Trees_din <= "00000000010100010101000001010101";
wait for Clk_period;
Addr <= "1010000000101";
Trees_din <= "00000000000010100101000001010101";
wait for Clk_period;
Addr <= "1010000000110";
Trees_din <= "00000001000000000100010000010000";
wait for Clk_period;
Addr <= "1010000000111";
Trees_din <= "00000110000000000000011000001000";
wait for Clk_period;
Addr <= "1010000001000";
Trees_din <= "00000001000000000010010000000100";
wait for Clk_period;
Addr <= "1010000001001";
Trees_din <= "00000000010111000101000001010101";
wait for Clk_period;
Addr <= "1010000001010";
Trees_din <= "00000000000101000101000001010101";
wait for Clk_period;
Addr <= "1010000001011";
Trees_din <= "00000111000000000010000100000100";
wait for Clk_period;
Addr <= "1010000001100";
Trees_din <= "00000000010011100101000001010101";
wait for Clk_period;
Addr <= "1010000001101";
Trees_din <= "00000000001110010101000001010101";
wait for Clk_period;
Addr <= "1010000001110";
Trees_din <= "00000001000000000010111000001000";
wait for Clk_period;
Addr <= "1010000001111";
Trees_din <= "00000100000000000100001100000100";
wait for Clk_period;
Addr <= "1010000010000";
Trees_din <= "00000000001001110101000001010101";
wait for Clk_period;
Addr <= "1010000010001";
Trees_din <= "00000000001110110101000001010101";
wait for Clk_period;
Addr <= "1010000010010";
Trees_din <= "00000000000000000010000000000100";
wait for Clk_period;
Addr <= "1010000010011";
Trees_din <= "00000000010101100101000001010101";
wait for Clk_period;
Addr <= "1010000010100";
Trees_din <= "00000000010011010101000001010101";
wait for Clk_period;



----------tree 40-------------------

Addr <= "1010000010101";
Trees_din <= "00000011000000000010011110000000";
wait for Clk_period;
Addr <= "1010000010110";
Trees_din <= "00000100000000000001000101000000";
wait for Clk_period;
Addr <= "1010000010111";
Trees_din <= "00000101000000000010010000100000";
wait for Clk_period;
Addr <= "1010000011000";
Trees_din <= "00000100000000000100010100010000";
wait for Clk_period;
Addr <= "1010000011001";
Trees_din <= "00000011000000000100011000001000";
wait for Clk_period;
Addr <= "1010000011010";
Trees_din <= "00000001000000000000010100000100";
wait for Clk_period;
Addr <= "1010000011011";
Trees_din <= "00000000001110010101001001010001";
wait for Clk_period;
Addr <= "1010000011100";
Trees_din <= "00000000001010100101001001010001";
wait for Clk_period;
Addr <= "1010000011101";
Trees_din <= "00000111000000000001101100000100";
wait for Clk_period;
Addr <= "1010000011110";
Trees_din <= "00000000010101010101001001010001";
wait for Clk_period;
Addr <= "1010000011111";
Trees_din <= "00000000001001100101001001010001";
wait for Clk_period;
Addr <= "1010000100000";
Trees_din <= "00000101000000000011001100001000";
wait for Clk_period;
Addr <= "1010000100001";
Trees_din <= "00000100000000000001101100000100";
wait for Clk_period;
Addr <= "1010000100010";
Trees_din <= "00000000000011010101001001010001";
wait for Clk_period;
Addr <= "1010000100011";
Trees_din <= "00000000000011000101001001010001";
wait for Clk_period;
Addr <= "1010000100100";
Trees_din <= "00000110000000000010110000000100";
wait for Clk_period;
Addr <= "1010000100101";
Trees_din <= "00000000000100100101001001010001";
wait for Clk_period;
Addr <= "1010000100110";
Trees_din <= "00000000000110100101001001010001";
wait for Clk_period;
Addr <= "1010000100111";
Trees_din <= "00000000000000000000100000010000";
wait for Clk_period;
Addr <= "1010000101000";
Trees_din <= "00000011000000000101101000001000";
wait for Clk_period;
Addr <= "1010000101001";
Trees_din <= "00000100000000000101001100000100";
wait for Clk_period;
Addr <= "1010000101010";
Trees_din <= "00000000001001000101001001010001";
wait for Clk_period;
Addr <= "1010000101011";
Trees_din <= "00000000010110010101001001010001";
wait for Clk_period;
Addr <= "1010000101100";
Trees_din <= "00000110000000000001010100000100";
wait for Clk_period;
Addr <= "1010000101101";
Trees_din <= "00000000001110000101001001010001";
wait for Clk_period;
Addr <= "1010000101110";
Trees_din <= "00000000000101110101001001010001";
wait for Clk_period;
Addr <= "1010000101111";
Trees_din <= "00000011000000000100100000001000";
wait for Clk_period;
Addr <= "1010000110000";
Trees_din <= "00000010000000000010010000000100";
wait for Clk_period;
Addr <= "1010000110001";
Trees_din <= "00000000001000010101001001010001";
wait for Clk_period;
Addr <= "1010000110010";
Trees_din <= "00000000000010100101001001010001";
wait for Clk_period;
Addr <= "1010000110011";
Trees_din <= "00000101000000000011000000000100";
wait for Clk_period;
Addr <= "1010000110100";
Trees_din <= "00000000001111010101001001010001";
wait for Clk_period;
Addr <= "1010000110101";
Trees_din <= "00000000010000000101001001010001";
wait for Clk_period;
Addr <= "1010000110110";
Trees_din <= "00000100000000000010011000100000";
wait for Clk_period;
Addr <= "1010000110111";
Trees_din <= "00000000000000000001101000010000";
wait for Clk_period;
Addr <= "1010000111000";
Trees_din <= "00000010000000000011101100001000";
wait for Clk_period;
Addr <= "1010000111001";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "1010000111010";
Trees_din <= "00000000000001110101001001010001";
wait for Clk_period;
Addr <= "1010000111011";
Trees_din <= "00000000000000000101001001010001";
wait for Clk_period;
Addr <= "1010000111100";
Trees_din <= "00000111000000000000110100000100";
wait for Clk_period;
Addr <= "1010000111101";
Trees_din <= "00000000001100000101001001010001";
wait for Clk_period;
Addr <= "1010000111110";
Trees_din <= "00000000010000000101001001010001";
wait for Clk_period;
Addr <= "1010000111111";
Trees_din <= "00000001000000000011001000001000";
wait for Clk_period;
Addr <= "1010001000000";
Trees_din <= "00000100000000000010010000000100";
wait for Clk_period;
Addr <= "1010001000001";
Trees_din <= "00000000000100110101001001010001";
wait for Clk_period;
Addr <= "1010001000010";
Trees_din <= "00000000000001110101001001010001";
wait for Clk_period;
Addr <= "1010001000011";
Trees_din <= "00000110000000000101000100000100";
wait for Clk_period;
Addr <= "1010001000100";
Trees_din <= "00000000000011110101001001010001";
wait for Clk_period;
Addr <= "1010001000101";
Trees_din <= "00000000000110100101001001010001";
wait for Clk_period;
Addr <= "1010001000110";
Trees_din <= "00000011000000000101110100010000";
wait for Clk_period;
Addr <= "1010001000111";
Trees_din <= "00000111000000000001101000001000";
wait for Clk_period;
Addr <= "1010001001000";
Trees_din <= "00000111000000000000101000000100";
wait for Clk_period;
Addr <= "1010001001001";
Trees_din <= "00000000011000010101001001010001";
wait for Clk_period;
Addr <= "1010001001010";
Trees_din <= "00000000010100100101001001010001";
wait for Clk_period;
Addr <= "1010001001011";
Trees_din <= "00000101000000000011101100000100";
wait for Clk_period;
Addr <= "1010001001100";
Trees_din <= "00000000000001010101001001010001";
wait for Clk_period;
Addr <= "1010001001101";
Trees_din <= "00000000000111110101001001010001";
wait for Clk_period;
Addr <= "1010001001110";
Trees_din <= "00000011000000000110001100001000";
wait for Clk_period;
Addr <= "1010001001111";
Trees_din <= "00000010000000000011101000000100";
wait for Clk_period;
Addr <= "1010001010000";
Trees_din <= "00000000011001000101001001010001";
wait for Clk_period;
Addr <= "1010001010001";
Trees_din <= "00000000010000110101001001010001";
wait for Clk_period;
Addr <= "1010001010010";
Trees_din <= "00000000000000000101011100000100";
wait for Clk_period;
Addr <= "1010001010011";
Trees_din <= "00000000000010010101001001010001";
wait for Clk_period;
Addr <= "1010001010100";
Trees_din <= "00000000000100110101001001010001";
wait for Clk_period;
Addr <= "1010001010101";
Trees_din <= "00000011000000000101001101000000";
wait for Clk_period;
Addr <= "1010001010110";
Trees_din <= "00000011000000000010011000100000";
wait for Clk_period;
Addr <= "1010001010111";
Trees_din <= "00000100000000000001001100010000";
wait for Clk_period;
Addr <= "1010001011000";
Trees_din <= "00000010000000000001010000001000";
wait for Clk_period;
Addr <= "1010001011001";
Trees_din <= "00000000000000000101111000000100";
wait for Clk_period;
Addr <= "1010001011010";
Trees_din <= "00000000010111110101001001010001";
wait for Clk_period;
Addr <= "1010001011011";
Trees_din <= "00000000000000000101001001010001";
wait for Clk_period;
Addr <= "1010001011100";
Trees_din <= "00000101000000000001001000000100";
wait for Clk_period;
Addr <= "1010001011101";
Trees_din <= "00000000001010000101001001010001";
wait for Clk_period;
Addr <= "1010001011110";
Trees_din <= "00000000011000000101001001010001";
wait for Clk_period;
Addr <= "1010001011111";
Trees_din <= "00000001000000000000101000001000";
wait for Clk_period;
Addr <= "1010001100000";
Trees_din <= "00000001000000000001100100000100";
wait for Clk_period;
Addr <= "1010001100001";
Trees_din <= "00000000001111100101001001010001";
wait for Clk_period;
Addr <= "1010001100010";
Trees_din <= "00000000000010010101001001010001";
wait for Clk_period;
Addr <= "1010001100011";
Trees_din <= "00000010000000000001111000000100";
wait for Clk_period;
Addr <= "1010001100100";
Trees_din <= "00000000010101110101001001010001";
wait for Clk_period;
Addr <= "1010001100101";
Trees_din <= "00000000000100110101001001010001";
wait for Clk_period;
Addr <= "1010001100110";
Trees_din <= "00000100000000000110001100010000";
wait for Clk_period;
Addr <= "1010001100111";
Trees_din <= "00000001000000000101011100001000";
wait for Clk_period;
Addr <= "1010001101000";
Trees_din <= "00000111000000000010111000000100";
wait for Clk_period;
Addr <= "1010001101001";
Trees_din <= "00000000000110110101001001010001";
wait for Clk_period;
Addr <= "1010001101010";
Trees_din <= "00000000010111100101001001010001";
wait for Clk_period;
Addr <= "1010001101011";
Trees_din <= "00000110000000000010100000000100";
wait for Clk_period;
Addr <= "1010001101100";
Trees_din <= "00000000001101100101001001010001";
wait for Clk_period;
Addr <= "1010001101101";
Trees_din <= "00000000010011010101001001010001";
wait for Clk_period;
Addr <= "1010001101110";
Trees_din <= "00000011000000000101001000001000";
wait for Clk_period;
Addr <= "1010001101111";
Trees_din <= "00000010000000000011101100000100";
wait for Clk_period;
Addr <= "1010001110000";
Trees_din <= "00000000000100110101001001010001";
wait for Clk_period;
Addr <= "1010001110001";
Trees_din <= "00000000000110010101001001010001";
wait for Clk_period;
Addr <= "1010001110010";
Trees_din <= "00000101000000000101011000000100";
wait for Clk_period;
Addr <= "1010001110011";
Trees_din <= "00000000010010100101001001010001";
wait for Clk_period;
Addr <= "1010001110100";
Trees_din <= "00000000000011010101001001010001";
wait for Clk_period;
Addr <= "1010001110101";
Trees_din <= "00000101000000000101010000100000";
wait for Clk_period;
Addr <= "1010001110110";
Trees_din <= "00000001000000000011000100010000";
wait for Clk_period;
Addr <= "1010001110111";
Trees_din <= "00000111000000000010000100001000";
wait for Clk_period;
Addr <= "1010001111000";
Trees_din <= "00000000000000000001001100000100";
wait for Clk_period;
Addr <= "1010001111001";
Trees_din <= "00000000010110010101001001010001";
wait for Clk_period;
Addr <= "1010001111010";
Trees_din <= "00000000000010010101001001010001";
wait for Clk_period;
Addr <= "1010001111011";
Trees_din <= "00000010000000000000000000000100";
wait for Clk_period;
Addr <= "1010001111100";
Trees_din <= "00000000001101000101001001010001";
wait for Clk_period;
Addr <= "1010001111101";
Trees_din <= "00000000001100110101001001010001";
wait for Clk_period;
Addr <= "1010001111110";
Trees_din <= "00000111000000000101001000001000";
wait for Clk_period;
Addr <= "1010001111111";
Trees_din <= "00000100000000000101011100000100";
wait for Clk_period;
Addr <= "1010010000000";
Trees_din <= "00000000000101010101001001010001";
wait for Clk_period;
Addr <= "1010010000001";
Trees_din <= "00000000001101110101001001010001";
wait for Clk_period;
Addr <= "1010010000010";
Trees_din <= "00000101000000000011011000000100";
wait for Clk_period;
Addr <= "1010010000011";
Trees_din <= "00000000010110100101001001010001";
wait for Clk_period;
Addr <= "1010010000100";
Trees_din <= "00000000000000010101001001010001";
wait for Clk_period;
Addr <= "1010010000101";
Trees_din <= "00000101000000000101000000010000";
wait for Clk_period;
Addr <= "1010010000110";
Trees_din <= "00000101000000000001100100001000";
wait for Clk_period;
Addr <= "1010010000111";
Trees_din <= "00000010000000000001000000000100";
wait for Clk_period;
Addr <= "1010010001000";
Trees_din <= "00000000000011000101001001010001";
wait for Clk_period;
Addr <= "1010010001001";
Trees_din <= "00000000000010100101001001010001";
wait for Clk_period;
Addr <= "1010010001010";
Trees_din <= "00000111000000000010111000000100";
wait for Clk_period;
Addr <= "1010010001011";
Trees_din <= "00000000010110010101001001010001";
wait for Clk_period;
Addr <= "1010010001100";
Trees_din <= "00000000001101010101001001010001";
wait for Clk_period;
Addr <= "1010010001101";
Trees_din <= "00000001000000000010011100001000";
wait for Clk_period;
Addr <= "1010010001110";
Trees_din <= "00000101000000000101100000000100";
wait for Clk_period;
Addr <= "1010010001111";
Trees_din <= "00000000010100110101001001010001";
wait for Clk_period;
Addr <= "1010010010000";
Trees_din <= "00000000010101000101001001010001";
wait for Clk_period;
Addr <= "1010010010001";
Trees_din <= "00000010000000000101100100000100";
wait for Clk_period;
Addr <= "1010010010010";
Trees_din <= "00000000000100010101001001010001";
wait for Clk_period;
Addr <= "1010010010011";
Trees_din <= "00000000001100000101001001010001";
wait for Clk_period;



----------tree 41-------------------

Addr <= "1010010010100";
Trees_din <= "00000010000000000100001110000000";
wait for Clk_period;
Addr <= "1010010010101";
Trees_din <= "00000110000000000101011001000000";
wait for Clk_period;
Addr <= "1010010010110";
Trees_din <= "00000000000000000101000000100000";
wait for Clk_period;
Addr <= "1010010010111";
Trees_din <= "00000010000000000010101000010000";
wait for Clk_period;
Addr <= "1010010011000";
Trees_din <= "00000110000000000100101100001000";
wait for Clk_period;
Addr <= "1010010011001";
Trees_din <= "00000000000000000000010000000100";
wait for Clk_period;
Addr <= "1010010011010";
Trees_din <= "00000000000100100101010001001101";
wait for Clk_period;
Addr <= "1010010011011";
Trees_din <= "00000000010000010101010001001101";
wait for Clk_period;
Addr <= "1010010011100";
Trees_din <= "00000000000000000100101100000100";
wait for Clk_period;
Addr <= "1010010011101";
Trees_din <= "00000000001111000101010001001101";
wait for Clk_period;
Addr <= "1010010011110";
Trees_din <= "00000000011001000101010001001101";
wait for Clk_period;
Addr <= "1010010011111";
Trees_din <= "00000010000000000010011000001000";
wait for Clk_period;
Addr <= "1010010100000";
Trees_din <= "00000011000000000010010000000100";
wait for Clk_period;
Addr <= "1010010100001";
Trees_din <= "00000000010001100101010001001101";
wait for Clk_period;
Addr <= "1010010100010";
Trees_din <= "00000000010011010101010001001101";
wait for Clk_period;
Addr <= "1010010100011";
Trees_din <= "00000010000000000000100000000100";
wait for Clk_period;
Addr <= "1010010100100";
Trees_din <= "00000000000101010101010001001101";
wait for Clk_period;
Addr <= "1010010100101";
Trees_din <= "00000000000111010101010001001101";
wait for Clk_period;
Addr <= "1010010100110";
Trees_din <= "00000101000000000100111000010000";
wait for Clk_period;
Addr <= "1010010100111";
Trees_din <= "00000101000000000000100100001000";
wait for Clk_period;
Addr <= "1010010101000";
Trees_din <= "00000001000000000100010000000100";
wait for Clk_period;
Addr <= "1010010101001";
Trees_din <= "00000000010110010101010001001101";
wait for Clk_period;
Addr <= "1010010101010";
Trees_din <= "00000000010101000101010001001101";
wait for Clk_period;
Addr <= "1010010101011";
Trees_din <= "00000111000000000011010000000100";
wait for Clk_period;
Addr <= "1010010101100";
Trees_din <= "00000000001011110101010001001101";
wait for Clk_period;
Addr <= "1010010101101";
Trees_din <= "00000000010001100101010001001101";
wait for Clk_period;
Addr <= "1010010101110";
Trees_din <= "00000110000000000101011100001000";
wait for Clk_period;
Addr <= "1010010101111";
Trees_din <= "00000111000000000110000000000100";
wait for Clk_period;
Addr <= "1010010110000";
Trees_din <= "00000000010001110101010001001101";
wait for Clk_period;
Addr <= "1010010110001";
Trees_din <= "00000000001011100101010001001101";
wait for Clk_period;
Addr <= "1010010110010";
Trees_din <= "00000101000000000101010000000100";
wait for Clk_period;
Addr <= "1010010110011";
Trees_din <= "00000000010010100101010001001101";
wait for Clk_period;
Addr <= "1010010110100";
Trees_din <= "00000000010001110101010001001101";
wait for Clk_period;
Addr <= "1010010110101";
Trees_din <= "00000011000000000010101000100000";
wait for Clk_period;
Addr <= "1010010110110";
Trees_din <= "00000000000000000110000000010000";
wait for Clk_period;
Addr <= "1010010110111";
Trees_din <= "00000011000000000010101000001000";
wait for Clk_period;
Addr <= "1010010111000";
Trees_din <= "00000001000000000011101000000100";
wait for Clk_period;
Addr <= "1010010111001";
Trees_din <= "00000000001010100101010001001101";
wait for Clk_period;
Addr <= "1010010111010";
Trees_din <= "00000000000011110101010001001101";
wait for Clk_period;
Addr <= "1010010111011";
Trees_din <= "00000100000000000001010000000100";
wait for Clk_period;
Addr <= "1010010111100";
Trees_din <= "00000000000111100101010001001101";
wait for Clk_period;
Addr <= "1010010111101";
Trees_din <= "00000000001010110101010001001101";
wait for Clk_period;
Addr <= "1010010111110";
Trees_din <= "00000101000000000101001100001000";
wait for Clk_period;
Addr <= "1010010111111";
Trees_din <= "00000011000000000101100000000100";
wait for Clk_period;
Addr <= "1010011000000";
Trees_din <= "00000000000110010101010001001101";
wait for Clk_period;
Addr <= "1010011000001";
Trees_din <= "00000000001000110101010001001101";
wait for Clk_period;
Addr <= "1010011000010";
Trees_din <= "00000011000000000011101100000100";
wait for Clk_period;
Addr <= "1010011000011";
Trees_din <= "00000000010101000101010001001101";
wait for Clk_period;
Addr <= "1010011000100";
Trees_din <= "00000000001010010101010001001101";
wait for Clk_period;
Addr <= "1010011000101";
Trees_din <= "00000100000000000100011100010000";
wait for Clk_period;
Addr <= "1010011000110";
Trees_din <= "00000001000000000100000000001000";
wait for Clk_period;
Addr <= "1010011000111";
Trees_din <= "00000101000000000110000000000100";
wait for Clk_period;
Addr <= "1010011001000";
Trees_din <= "00000000000111100101010001001101";
wait for Clk_period;
Addr <= "1010011001001";
Trees_din <= "00000000000111000101010001001101";
wait for Clk_period;
Addr <= "1010011001010";
Trees_din <= "00000001000000000011000000000100";
wait for Clk_period;
Addr <= "1010011001011";
Trees_din <= "00000000001001010101010001001101";
wait for Clk_period;
Addr <= "1010011001100";
Trees_din <= "00000000001010110101010001001101";
wait for Clk_period;
Addr <= "1010011001101";
Trees_din <= "00000001000000000000101000001000";
wait for Clk_period;
Addr <= "1010011001110";
Trees_din <= "00000100000000000000010000000100";
wait for Clk_period;
Addr <= "1010011001111";
Trees_din <= "00000000000001110101010001001101";
wait for Clk_period;
Addr <= "1010011010000";
Trees_din <= "00000000000000010101010001001101";
wait for Clk_period;
Addr <= "1010011010001";
Trees_din <= "00000111000000000010111100000100";
wait for Clk_period;
Addr <= "1010011010010";
Trees_din <= "00000000010010010101010001001101";
wait for Clk_period;
Addr <= "1010011010011";
Trees_din <= "00000000001010010101010001001101";
wait for Clk_period;
Addr <= "1010011010100";
Trees_din <= "00000111000000000011000001000000";
wait for Clk_period;
Addr <= "1010011010101";
Trees_din <= "00000001000000000000011000100000";
wait for Clk_period;
Addr <= "1010011010110";
Trees_din <= "00000111000000000001001000010000";
wait for Clk_period;
Addr <= "1010011010111";
Trees_din <= "00000011000000000101010000001000";
wait for Clk_period;
Addr <= "1010011011000";
Trees_din <= "00000111000000000110000100000100";
wait for Clk_period;
Addr <= "1010011011001";
Trees_din <= "00000000010100110101010001001101";
wait for Clk_period;
Addr <= "1010011011010";
Trees_din <= "00000000010100100101010001001101";
wait for Clk_period;
Addr <= "1010011011011";
Trees_din <= "00000101000000000001101100000100";
wait for Clk_period;
Addr <= "1010011011100";
Trees_din <= "00000000000011000101010001001101";
wait for Clk_period;
Addr <= "1010011011101";
Trees_din <= "00000000000111100101010001001101";
wait for Clk_period;
Addr <= "1010011011110";
Trees_din <= "00000111000000000000011100001000";
wait for Clk_period;
Addr <= "1010011011111";
Trees_din <= "00000100000000000010101000000100";
wait for Clk_period;
Addr <= "1010011100000";
Trees_din <= "00000000001000110101010001001101";
wait for Clk_period;
Addr <= "1010011100001";
Trees_din <= "00000000001100000101010001001101";
wait for Clk_period;
Addr <= "1010011100010";
Trees_din <= "00000101000000000101101100000100";
wait for Clk_period;
Addr <= "1010011100011";
Trees_din <= "00000000010000100101010001001101";
wait for Clk_period;
Addr <= "1010011100100";
Trees_din <= "00000000001001010101010001001101";
wait for Clk_period;
Addr <= "1010011100101";
Trees_din <= "00000000000000000011110000010000";
wait for Clk_period;
Addr <= "1010011100110";
Trees_din <= "00000111000000000011001100001000";
wait for Clk_period;
Addr <= "1010011100111";
Trees_din <= "00000110000000000100011100000100";
wait for Clk_period;
Addr <= "1010011101000";
Trees_din <= "00000000001001100101010001001101";
wait for Clk_period;
Addr <= "1010011101001";
Trees_din <= "00000000001000010101010001001101";
wait for Clk_period;
Addr <= "1010011101010";
Trees_din <= "00000100000000000100011100000100";
wait for Clk_period;
Addr <= "1010011101011";
Trees_din <= "00000000011000110101010001001101";
wait for Clk_period;
Addr <= "1010011101100";
Trees_din <= "00000000000110110101010001001101";
wait for Clk_period;
Addr <= "1010011101101";
Trees_din <= "00000100000000000010001100001000";
wait for Clk_period;
Addr <= "1010011101110";
Trees_din <= "00000101000000000101001000000100";
wait for Clk_period;
Addr <= "1010011101111";
Trees_din <= "00000000011000010101010001001101";
wait for Clk_period;
Addr <= "1010011110000";
Trees_din <= "00000000010001010101010001001101";
wait for Clk_period;
Addr <= "1010011110001";
Trees_din <= "00000100000000000011111000000100";
wait for Clk_period;
Addr <= "1010011110010";
Trees_din <= "00000000010010010101010001001101";
wait for Clk_period;
Addr <= "1010011110011";
Trees_din <= "00000000001100100101010001001101";
wait for Clk_period;
Addr <= "1010011110100";
Trees_din <= "00000111000000000101010000100000";
wait for Clk_period;
Addr <= "1010011110101";
Trees_din <= "00000100000000000110001000010000";
wait for Clk_period;
Addr <= "1010011110110";
Trees_din <= "00000100000000000011110100001000";
wait for Clk_period;
Addr <= "1010011110111";
Trees_din <= "00000010000000000000001000000100";
wait for Clk_period;
Addr <= "1010011111000";
Trees_din <= "00000000000111010101010001001101";
wait for Clk_period;
Addr <= "1010011111001";
Trees_din <= "00000000000000010101010001001101";
wait for Clk_period;
Addr <= "1010011111010";
Trees_din <= "00000000000000000001101100000100";
wait for Clk_period;
Addr <= "1010011111011";
Trees_din <= "00000000000001100101010001001101";
wait for Clk_period;
Addr <= "1010011111100";
Trees_din <= "00000000000001000101010001001101";
wait for Clk_period;
Addr <= "1010011111101";
Trees_din <= "00000010000000000000100000001000";
wait for Clk_period;
Addr <= "1010011111110";
Trees_din <= "00000000000000000100000000000100";
wait for Clk_period;
Addr <= "1010011111111";
Trees_din <= "00000000010110100101010001001101";
wait for Clk_period;
Addr <= "1010100000000";
Trees_din <= "00000000010010000101010001001101";
wait for Clk_period;
Addr <= "1010100000001";
Trees_din <= "00000000000000000000101000000100";
wait for Clk_period;
Addr <= "1010100000010";
Trees_din <= "00000000001001010101010001001101";
wait for Clk_period;
Addr <= "1010100000011";
Trees_din <= "00000000010000010101010001001101";
wait for Clk_period;
Addr <= "1010100000100";
Trees_din <= "00000111000000000000010100010000";
wait for Clk_period;
Addr <= "1010100000101";
Trees_din <= "00000011000000000101001100001000";
wait for Clk_period;
Addr <= "1010100000110";
Trees_din <= "00000000000000000110001100000100";
wait for Clk_period;
Addr <= "1010100000111";
Trees_din <= "00000000010110110101010001001101";
wait for Clk_period;
Addr <= "1010100001000";
Trees_din <= "00000000001101010101010001001101";
wait for Clk_period;
Addr <= "1010100001001";
Trees_din <= "00000100000000000101111000000100";
wait for Clk_period;
Addr <= "1010100001010";
Trees_din <= "00000000001100110101010001001101";
wait for Clk_period;
Addr <= "1010100001011";
Trees_din <= "00000000011000010101010001001101";
wait for Clk_period;
Addr <= "1010100001100";
Trees_din <= "00000001000000000001000000001000";
wait for Clk_period;
Addr <= "1010100001101";
Trees_din <= "00000100000000000101010000000100";
wait for Clk_period;
Addr <= "1010100001110";
Trees_din <= "00000000010110100101010001001101";
wait for Clk_period;
Addr <= "1010100001111";
Trees_din <= "00000000010010000101010001001101";
wait for Clk_period;
Addr <= "1010100010000";
Trees_din <= "00000001000000000010110000000100";
wait for Clk_period;
Addr <= "1010100010001";
Trees_din <= "00000000000010000101010001001101";
wait for Clk_period;
Addr <= "1010100010010";
Trees_din <= "00000000000111000101010001001101";
wait for Clk_period;



----------tree 42-------------------

Addr <= "1010100010011";
Trees_din <= "00000101000000000010011110000000";
wait for Clk_period;
Addr <= "1010100010100";
Trees_din <= "00000010000000000000010101000000";
wait for Clk_period;
Addr <= "1010100010101";
Trees_din <= "00000011000000000101010100100000";
wait for Clk_period;
Addr <= "1010100010110";
Trees_din <= "00000111000000000011000000010000";
wait for Clk_period;
Addr <= "1010100010111";
Trees_din <= "00000001000000000000000100001000";
wait for Clk_period;
Addr <= "1010100011000";
Trees_din <= "00000111000000000001011100000100";
wait for Clk_period;
Addr <= "1010100011001";
Trees_din <= "00000000000100100101011001001001";
wait for Clk_period;
Addr <= "1010100011010";
Trees_din <= "00000000000000000101011001001001";
wait for Clk_period;
Addr <= "1010100011011";
Trees_din <= "00000000000000000101011000000100";
wait for Clk_period;
Addr <= "1010100011100";
Trees_din <= "00000000010101000101011001001001";
wait for Clk_period;
Addr <= "1010100011101";
Trees_din <= "00000000000011010101011001001001";
wait for Clk_period;
Addr <= "1010100011110";
Trees_din <= "00000101000000000000100100001000";
wait for Clk_period;
Addr <= "1010100011111";
Trees_din <= "00000111000000000101100100000100";
wait for Clk_period;
Addr <= "1010100100000";
Trees_din <= "00000000010001010101011001001001";
wait for Clk_period;
Addr <= "1010100100001";
Trees_din <= "00000000001111000101011001001001";
wait for Clk_period;
Addr <= "1010100100010";
Trees_din <= "00000110000000000100111100000100";
wait for Clk_period;
Addr <= "1010100100011";
Trees_din <= "00000000000001110101011001001001";
wait for Clk_period;
Addr <= "1010100100100";
Trees_din <= "00000000001001000101011001001001";
wait for Clk_period;
Addr <= "1010100100101";
Trees_din <= "00000001000000000101001000010000";
wait for Clk_period;
Addr <= "1010100100110";
Trees_din <= "00000011000000000011101000001000";
wait for Clk_period;
Addr <= "1010100100111";
Trees_din <= "00000000000000000101011000000100";
wait for Clk_period;
Addr <= "1010100101000";
Trees_din <= "00000000001100100101011001001001";
wait for Clk_period;
Addr <= "1010100101001";
Trees_din <= "00000000001111100101011001001001";
wait for Clk_period;
Addr <= "1010100101010";
Trees_din <= "00000100000000000011100100000100";
wait for Clk_period;
Addr <= "1010100101011";
Trees_din <= "00000000010100100101011001001001";
wait for Clk_period;
Addr <= "1010100101100";
Trees_din <= "00000000010101110101011001001001";
wait for Clk_period;
Addr <= "1010100101101";
Trees_din <= "00000101000000000100111000001000";
wait for Clk_period;
Addr <= "1010100101110";
Trees_din <= "00000101000000000010011100000100";
wait for Clk_period;
Addr <= "1010100101111";
Trees_din <= "00000000010111010101011001001001";
wait for Clk_period;
Addr <= "1010100110000";
Trees_din <= "00000000010011100101011001001001";
wait for Clk_period;
Addr <= "1010100110001";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "1010100110010";
Trees_din <= "00000000010110100101011001001001";
wait for Clk_period;
Addr <= "1010100110011";
Trees_din <= "00000000001101000101011001001001";
wait for Clk_period;
Addr <= "1010100110100";
Trees_din <= "00000100000000000100001100100000";
wait for Clk_period;
Addr <= "1010100110101";
Trees_din <= "00000111000000000000100100010000";
wait for Clk_period;
Addr <= "1010100110110";
Trees_din <= "00000001000000000001000100001000";
wait for Clk_period;
Addr <= "1010100110111";
Trees_din <= "00000110000000000001111000000100";
wait for Clk_period;
Addr <= "1010100111000";
Trees_din <= "00000000000100010101011001001001";
wait for Clk_period;
Addr <= "1010100111001";
Trees_din <= "00000000001100010101011001001001";
wait for Clk_period;
Addr <= "1010100111010";
Trees_din <= "00000000000000000101100100000100";
wait for Clk_period;
Addr <= "1010100111011";
Trees_din <= "00000000010000010101011001001001";
wait for Clk_period;
Addr <= "1010100111100";
Trees_din <= "00000000010101110101011001001001";
wait for Clk_period;
Addr <= "1010100111101";
Trees_din <= "00000011000000000011000100001000";
wait for Clk_period;
Addr <= "1010100111110";
Trees_din <= "00000100000000000011011000000100";
wait for Clk_period;
Addr <= "1010100111111";
Trees_din <= "00000000001001010101011001001001";
wait for Clk_period;
Addr <= "1010101000000";
Trees_din <= "00000000011000010101011001001001";
wait for Clk_period;
Addr <= "1010101000001";
Trees_din <= "00000110000000000100000100000100";
wait for Clk_period;
Addr <= "1010101000010";
Trees_din <= "00000000010100000101011001001001";
wait for Clk_period;
Addr <= "1010101000011";
Trees_din <= "00000000000111110101011001001001";
wait for Clk_period;
Addr <= "1010101000100";
Trees_din <= "00000011000000000110001100010000";
wait for Clk_period;
Addr <= "1010101000101";
Trees_din <= "00000100000000000011011100001000";
wait for Clk_period;
Addr <= "1010101000110";
Trees_din <= "00000110000000000010111100000100";
wait for Clk_period;
Addr <= "1010101000111";
Trees_din <= "00000000010001110101011001001001";
wait for Clk_period;
Addr <= "1010101001000";
Trees_din <= "00000000010001110101011001001001";
wait for Clk_period;
Addr <= "1010101001001";
Trees_din <= "00000001000000000010010000000100";
wait for Clk_period;
Addr <= "1010101001010";
Trees_din <= "00000000000010000101011001001001";
wait for Clk_period;
Addr <= "1010101001011";
Trees_din <= "00000000000011100101011001001001";
wait for Clk_period;
Addr <= "1010101001100";
Trees_din <= "00000111000000000000001100001000";
wait for Clk_period;
Addr <= "1010101001101";
Trees_din <= "00000111000000000100000100000100";
wait for Clk_period;
Addr <= "1010101001110";
Trees_din <= "00000000010110000101011001001001";
wait for Clk_period;
Addr <= "1010101001111";
Trees_din <= "00000000011000110101011001001001";
wait for Clk_period;
Addr <= "1010101010000";
Trees_din <= "00000010000000000001111000000100";
wait for Clk_period;
Addr <= "1010101010001";
Trees_din <= "00000000010111000101011001001001";
wait for Clk_period;
Addr <= "1010101010010";
Trees_din <= "00000000000001110101011001001001";
wait for Clk_period;
Addr <= "1010101010011";
Trees_din <= "00000100000000000101010001000000";
wait for Clk_period;
Addr <= "1010101010100";
Trees_din <= "00000110000000000101001100100000";
wait for Clk_period;
Addr <= "1010101010101";
Trees_din <= "00000100000000000101100000010000";
wait for Clk_period;
Addr <= "1010101010110";
Trees_din <= "00000000000000000010011000001000";
wait for Clk_period;
Addr <= "1010101010111";
Trees_din <= "00000111000000000101011100000100";
wait for Clk_period;
Addr <= "1010101011000";
Trees_din <= "00000000001111000101011001001001";
wait for Clk_period;
Addr <= "1010101011001";
Trees_din <= "00000000010011100101011001001001";
wait for Clk_period;
Addr <= "1010101011010";
Trees_din <= "00000011000000000110010000000100";
wait for Clk_period;
Addr <= "1010101011011";
Trees_din <= "00000000011000100101011001001001";
wait for Clk_period;
Addr <= "1010101011100";
Trees_din <= "00000000010001110101011001001001";
wait for Clk_period;
Addr <= "1010101011101";
Trees_din <= "00000000000000000100001100001000";
wait for Clk_period;
Addr <= "1010101011110";
Trees_din <= "00000101000000000101011100000100";
wait for Clk_period;
Addr <= "1010101011111";
Trees_din <= "00000000000011100101011001001001";
wait for Clk_period;
Addr <= "1010101100000";
Trees_din <= "00000000000111110101011001001001";
wait for Clk_period;
Addr <= "1010101100001";
Trees_din <= "00000100000000000000101000000100";
wait for Clk_period;
Addr <= "1010101100010";
Trees_din <= "00000000000001000101011001001001";
wait for Clk_period;
Addr <= "1010101100011";
Trees_din <= "00000000001100100101011001001001";
wait for Clk_period;
Addr <= "1010101100100";
Trees_din <= "00000110000000000100010000010000";
wait for Clk_period;
Addr <= "1010101100101";
Trees_din <= "00000000000000000011100100001000";
wait for Clk_period;
Addr <= "1010101100110";
Trees_din <= "00000011000000000001010000000100";
wait for Clk_period;
Addr <= "1010101100111";
Trees_din <= "00000000000111100101011001001001";
wait for Clk_period;
Addr <= "1010101101000";
Trees_din <= "00000000011001000101011001001001";
wait for Clk_period;
Addr <= "1010101101001";
Trees_din <= "00000101000000000001101000000100";
wait for Clk_period;
Addr <= "1010101101010";
Trees_din <= "00000000001111000101011001001001";
wait for Clk_period;
Addr <= "1010101101011";
Trees_din <= "00000000010101010101011001001001";
wait for Clk_period;
Addr <= "1010101101100";
Trees_din <= "00000011000000000001001100001000";
wait for Clk_period;
Addr <= "1010101101101";
Trees_din <= "00000000000000000100001000000100";
wait for Clk_period;
Addr <= "1010101101110";
Trees_din <= "00000000000101110101011001001001";
wait for Clk_period;
Addr <= "1010101101111";
Trees_din <= "00000000010111000101011001001001";
wait for Clk_period;
Addr <= "1010101110000";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "1010101110001";
Trees_din <= "00000000010111000101011001001001";
wait for Clk_period;
Addr <= "1010101110010";
Trees_din <= "00000000001111100101011001001001";
wait for Clk_period;
Addr <= "1010101110011";
Trees_din <= "00000100000000000100101100100000";
wait for Clk_period;
Addr <= "1010101110100";
Trees_din <= "00000110000000000001001000010000";
wait for Clk_period;
Addr <= "1010101110101";
Trees_din <= "00000010000000000101110100001000";
wait for Clk_period;
Addr <= "1010101110110";
Trees_din <= "00000100000000000101010000000100";
wait for Clk_period;
Addr <= "1010101110111";
Trees_din <= "00000000010001110101011001001001";
wait for Clk_period;
Addr <= "1010101111000";
Trees_din <= "00000000010100010101011001001001";
wait for Clk_period;
Addr <= "1010101111001";
Trees_din <= "00000111000000000011111000000100";
wait for Clk_period;
Addr <= "1010101111010";
Trees_din <= "00000000000001000101011001001001";
wait for Clk_period;
Addr <= "1010101111011";
Trees_din <= "00000000001100100101011001001001";
wait for Clk_period;
Addr <= "1010101111100";
Trees_din <= "00000000000000000011111100001000";
wait for Clk_period;
Addr <= "1010101111101";
Trees_din <= "00000011000000000011010100000100";
wait for Clk_period;
Addr <= "1010101111110";
Trees_din <= "00000000010000010101011001001001";
wait for Clk_period;
Addr <= "1010101111111";
Trees_din <= "00000000011000000101011001001001";
wait for Clk_period;
Addr <= "1010110000000";
Trees_din <= "00000100000000000010000100000100";
wait for Clk_period;
Addr <= "1010110000001";
Trees_din <= "00000000000111110101011001001001";
wait for Clk_period;
Addr <= "1010110000010";
Trees_din <= "00000000010001010101011001001001";
wait for Clk_period;
Addr <= "1010110000011";
Trees_din <= "00000010000000000001000100010000";
wait for Clk_period;
Addr <= "1010110000100";
Trees_din <= "00000111000000000001001100001000";
wait for Clk_period;
Addr <= "1010110000101";
Trees_din <= "00000001000000000011010100000100";
wait for Clk_period;
Addr <= "1010110000110";
Trees_din <= "00000000000100110101011001001001";
wait for Clk_period;
Addr <= "1010110000111";
Trees_din <= "00000000010111010101011001001001";
wait for Clk_period;
Addr <= "1010110001000";
Trees_din <= "00000001000000000000010100000100";
wait for Clk_period;
Addr <= "1010110001001";
Trees_din <= "00000000000100100101011001001001";
wait for Clk_period;
Addr <= "1010110001010";
Trees_din <= "00000000000000110101011001001001";
wait for Clk_period;
Addr <= "1010110001011";
Trees_din <= "00000011000000000010101000001000";
wait for Clk_period;
Addr <= "1010110001100";
Trees_din <= "00000001000000000101111100000100";
wait for Clk_period;
Addr <= "1010110001101";
Trees_din <= "00000000010011100101011001001001";
wait for Clk_period;
Addr <= "1010110001110";
Trees_din <= "00000000001011100101011001001001";
wait for Clk_period;
Addr <= "1010110001111";
Trees_din <= "00000100000000000011111000000100";
wait for Clk_period;
Addr <= "1010110010000";
Trees_din <= "00000000011000000101011001001001";
wait for Clk_period;
Addr <= "1010110010001";
Trees_din <= "00000000000101000101011001001001";
wait for Clk_period;



----------tree 43-------------------

Addr <= "1010110010010";
Trees_din <= "00000000000000000101101110000000";
wait for Clk_period;
Addr <= "1010110010011";
Trees_din <= "00000101000000000011010001000000";
wait for Clk_period;
Addr <= "1010110010100";
Trees_din <= "00000011000000000000000000100000";
wait for Clk_period;
Addr <= "1010110010101";
Trees_din <= "00000110000000000101110100010000";
wait for Clk_period;
Addr <= "1010110010110";
Trees_din <= "00000110000000000001101100001000";
wait for Clk_period;
Addr <= "1010110010111";
Trees_din <= "00000111000000000101001100000100";
wait for Clk_period;
Addr <= "1010110011000";
Trees_din <= "00000000010111010101100001000101";
wait for Clk_period;
Addr <= "1010110011001";
Trees_din <= "00000000010101100101100001000101";
wait for Clk_period;
Addr <= "1010110011010";
Trees_din <= "00000101000000000101101100000100";
wait for Clk_period;
Addr <= "1010110011011";
Trees_din <= "00000000010100000101100001000101";
wait for Clk_period;
Addr <= "1010110011100";
Trees_din <= "00000000011000000101100001000101";
wait for Clk_period;
Addr <= "1010110011101";
Trees_din <= "00000101000000000000001100001000";
wait for Clk_period;
Addr <= "1010110011110";
Trees_din <= "00000010000000000100111000000100";
wait for Clk_period;
Addr <= "1010110011111";
Trees_din <= "00000000000111010101100001000101";
wait for Clk_period;
Addr <= "1010110100000";
Trees_din <= "00000000000011100101100001000101";
wait for Clk_period;
Addr <= "1010110100001";
Trees_din <= "00000111000000000011101100000100";
wait for Clk_period;
Addr <= "1010110100010";
Trees_din <= "00000000011001000101100001000101";
wait for Clk_period;
Addr <= "1010110100011";
Trees_din <= "00000000010110000101100001000101";
wait for Clk_period;
Addr <= "1010110100100";
Trees_din <= "00000000000000000110010000010000";
wait for Clk_period;
Addr <= "1010110100101";
Trees_din <= "00000101000000000001111100001000";
wait for Clk_period;
Addr <= "1010110100110";
Trees_din <= "00000010000000000011001100000100";
wait for Clk_period;
Addr <= "1010110100111";
Trees_din <= "00000000000110000101100001000101";
wait for Clk_period;
Addr <= "1010110101000";
Trees_din <= "00000000001110100101100001000101";
wait for Clk_period;
Addr <= "1010110101001";
Trees_din <= "00000110000000000010001100000100";
wait for Clk_period;
Addr <= "1010110101010";
Trees_din <= "00000000010110010101100001000101";
wait for Clk_period;
Addr <= "1010110101011";
Trees_din <= "00000000001011010101100001000101";
wait for Clk_period;
Addr <= "1010110101100";
Trees_din <= "00000111000000000100100000001000";
wait for Clk_period;
Addr <= "1010110101101";
Trees_din <= "00000110000000000000000100000100";
wait for Clk_period;
Addr <= "1010110101110";
Trees_din <= "00000000010111010101100001000101";
wait for Clk_period;
Addr <= "1010110101111";
Trees_din <= "00000000000111100101100001000101";
wait for Clk_period;
Addr <= "1010110110000";
Trees_din <= "00000100000000000100111100000100";
wait for Clk_period;
Addr <= "1010110110001";
Trees_din <= "00000000010011100101100001000101";
wait for Clk_period;
Addr <= "1010110110010";
Trees_din <= "00000000011000110101100001000101";
wait for Clk_period;
Addr <= "1010110110011";
Trees_din <= "00000001000000000101101100100000";
wait for Clk_period;
Addr <= "1010110110100";
Trees_din <= "00000010000000000101000100010000";
wait for Clk_period;
Addr <= "1010110110101";
Trees_din <= "00000111000000000010010000001000";
wait for Clk_period;
Addr <= "1010110110110";
Trees_din <= "00000111000000000101011100000100";
wait for Clk_period;
Addr <= "1010110110111";
Trees_din <= "00000000000110000101100001000101";
wait for Clk_period;
Addr <= "1010110111000";
Trees_din <= "00000000001111110101100001000101";
wait for Clk_period;
Addr <= "1010110111001";
Trees_din <= "00000111000000000011001100000100";
wait for Clk_period;
Addr <= "1010110111010";
Trees_din <= "00000000001001100101100001000101";
wait for Clk_period;
Addr <= "1010110111011";
Trees_din <= "00000000000111010101100001000101";
wait for Clk_period;
Addr <= "1010110111100";
Trees_din <= "00000011000000000110000100001000";
wait for Clk_period;
Addr <= "1010110111101";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "1010110111110";
Trees_din <= "00000000001000010101100001000101";
wait for Clk_period;
Addr <= "1010110111111";
Trees_din <= "00000000000000010101100001000101";
wait for Clk_period;
Addr <= "1010111000000";
Trees_din <= "00000010000000000000001000000100";
wait for Clk_period;
Addr <= "1010111000001";
Trees_din <= "00000000001100010101100001000101";
wait for Clk_period;
Addr <= "1010111000010";
Trees_din <= "00000000000011010101100001000101";
wait for Clk_period;
Addr <= "1010111000011";
Trees_din <= "00000011000000000011010100010000";
wait for Clk_period;
Addr <= "1010111000100";
Trees_din <= "00000001000000000110000000001000";
wait for Clk_period;
Addr <= "1010111000101";
Trees_din <= "00000010000000000100001000000100";
wait for Clk_period;
Addr <= "1010111000110";
Trees_din <= "00000000001111100101100001000101";
wait for Clk_period;
Addr <= "1010111000111";
Trees_din <= "00000000000101010101100001000101";
wait for Clk_period;
Addr <= "1010111001000";
Trees_din <= "00000101000000000010001000000100";
wait for Clk_period;
Addr <= "1010111001001";
Trees_din <= "00000000010101010101100001000101";
wait for Clk_period;
Addr <= "1010111001010";
Trees_din <= "00000000000001000101100001000101";
wait for Clk_period;
Addr <= "1010111001011";
Trees_din <= "00000011000000000100101000001000";
wait for Clk_period;
Addr <= "1010111001100";
Trees_din <= "00000001000000000001110100000100";
wait for Clk_period;
Addr <= "1010111001101";
Trees_din <= "00000000001110100101100001000101";
wait for Clk_period;
Addr <= "1010111001110";
Trees_din <= "00000000010011010101100001000101";
wait for Clk_period;
Addr <= "1010111001111";
Trees_din <= "00000001000000000000000000000100";
wait for Clk_period;
Addr <= "1010111010000";
Trees_din <= "00000000000101010101100001000101";
wait for Clk_period;
Addr <= "1010111010001";
Trees_din <= "00000000010101110101100001000101";
wait for Clk_period;
Addr <= "1010111010010";
Trees_din <= "00000010000000000100000101000000";
wait for Clk_period;
Addr <= "1010111010011";
Trees_din <= "00000010000000000100001000100000";
wait for Clk_period;
Addr <= "1010111010100";
Trees_din <= "00000110000000000001010000010000";
wait for Clk_period;
Addr <= "1010111010101";
Trees_din <= "00000110000000000100110000001000";
wait for Clk_period;
Addr <= "1010111010110";
Trees_din <= "00000110000000000000000100000100";
wait for Clk_period;
Addr <= "1010111010111";
Trees_din <= "00000000000110010101100001000101";
wait for Clk_period;
Addr <= "1010111011000";
Trees_din <= "00000000000000110101100001000101";
wait for Clk_period;
Addr <= "1010111011001";
Trees_din <= "00000010000000000110000100000100";
wait for Clk_period;
Addr <= "1010111011010";
Trees_din <= "00000000010000000101100001000101";
wait for Clk_period;
Addr <= "1010111011011";
Trees_din <= "00000000000110110101100001000101";
wait for Clk_period;
Addr <= "1010111011100";
Trees_din <= "00000001000000000100011000001000";
wait for Clk_period;
Addr <= "1010111011101";
Trees_din <= "00000011000000000011001100000100";
wait for Clk_period;
Addr <= "1010111011110";
Trees_din <= "00000000001100110101100001000101";
wait for Clk_period;
Addr <= "1010111011111";
Trees_din <= "00000000010111000101100001000101";
wait for Clk_period;
Addr <= "1010111100000";
Trees_din <= "00000000000000000000001000000100";
wait for Clk_period;
Addr <= "1010111100001";
Trees_din <= "00000000001010110101100001000101";
wait for Clk_period;
Addr <= "1010111100010";
Trees_din <= "00000000000100000101100001000101";
wait for Clk_period;
Addr <= "1010111100011";
Trees_din <= "00000011000000000010000000010000";
wait for Clk_period;
Addr <= "1010111100100";
Trees_din <= "00000001000000000011001000001000";
wait for Clk_period;
Addr <= "1010111100101";
Trees_din <= "00000010000000000101001100000100";
wait for Clk_period;
Addr <= "1010111100110";
Trees_din <= "00000000010100010101100001000101";
wait for Clk_period;
Addr <= "1010111100111";
Trees_din <= "00000000001110100101100001000101";
wait for Clk_period;
Addr <= "1010111101000";
Trees_din <= "00000101000000000000110100000100";
wait for Clk_period;
Addr <= "1010111101001";
Trees_din <= "00000000000101100101100001000101";
wait for Clk_period;
Addr <= "1010111101010";
Trees_din <= "00000000001111010101100001000101";
wait for Clk_period;
Addr <= "1010111101011";
Trees_din <= "00000110000000000011001100001000";
wait for Clk_period;
Addr <= "1010111101100";
Trees_din <= "00000001000000000110000100000100";
wait for Clk_period;
Addr <= "1010111101101";
Trees_din <= "00000000010100010101100001000101";
wait for Clk_period;
Addr <= "1010111101110";
Trees_din <= "00000000010110100101100001000101";
wait for Clk_period;
Addr <= "1010111101111";
Trees_din <= "00000110000000000000001000000100";
wait for Clk_period;
Addr <= "1010111110000";
Trees_din <= "00000000001101010101100001000101";
wait for Clk_period;
Addr <= "1010111110001";
Trees_din <= "00000000000001100101100001000101";
wait for Clk_period;
Addr <= "1010111110010";
Trees_din <= "00000111000000000010001000100000";
wait for Clk_period;
Addr <= "1010111110011";
Trees_din <= "00000100000000000000011000010000";
wait for Clk_period;
Addr <= "1010111110100";
Trees_din <= "00000000000000000001110100001000";
wait for Clk_period;
Addr <= "1010111110101";
Trees_din <= "00000011000000000110000000000100";
wait for Clk_period;
Addr <= "1010111110110";
Trees_din <= "00000000000011010101100001000101";
wait for Clk_period;
Addr <= "1010111110111";
Trees_din <= "00000000011000100101100001000101";
wait for Clk_period;
Addr <= "1010111111000";
Trees_din <= "00000110000000000011111000000100";
wait for Clk_period;
Addr <= "1010111111001";
Trees_din <= "00000000001001000101100001000101";
wait for Clk_period;
Addr <= "1010111111010";
Trees_din <= "00000000000011010101100001000101";
wait for Clk_period;
Addr <= "1010111111011";
Trees_din <= "00000110000000000101000000001000";
wait for Clk_period;
Addr <= "1010111111100";
Trees_din <= "00000111000000000101001100000100";
wait for Clk_period;
Addr <= "1010111111101";
Trees_din <= "00000000001000010101100001000101";
wait for Clk_period;
Addr <= "1010111111110";
Trees_din <= "00000000001111100101100001000101";
wait for Clk_period;
Addr <= "1010111111111";
Trees_din <= "00000011000000000010111000000100";
wait for Clk_period;
Addr <= "1011000000000";
Trees_din <= "00000000000111100101100001000101";
wait for Clk_period;
Addr <= "1011000000001";
Trees_din <= "00000000011000100101100001000101";
wait for Clk_period;
Addr <= "1011000000010";
Trees_din <= "00000000000000000100100000010000";
wait for Clk_period;
Addr <= "1011000000011";
Trees_din <= "00000111000000000011001100001000";
wait for Clk_period;
Addr <= "1011000000100";
Trees_din <= "00000101000000000010001100000100";
wait for Clk_period;
Addr <= "1011000000101";
Trees_din <= "00000000010110110101100001000101";
wait for Clk_period;
Addr <= "1011000000110";
Trees_din <= "00000000000100000101100001000101";
wait for Clk_period;
Addr <= "1011000000111";
Trees_din <= "00000101000000000001100000000100";
wait for Clk_period;
Addr <= "1011000001000";
Trees_din <= "00000000000001110101100001000101";
wait for Clk_period;
Addr <= "1011000001001";
Trees_din <= "00000000011000100101100001000101";
wait for Clk_period;
Addr <= "1011000001010";
Trees_din <= "00000011000000000011001000001000";
wait for Clk_period;
Addr <= "1011000001011";
Trees_din <= "00000110000000000010011100000100";
wait for Clk_period;
Addr <= "1011000001100";
Trees_din <= "00000000001010110101100001000101";
wait for Clk_period;
Addr <= "1011000001101";
Trees_din <= "00000000000111010101100001000101";
wait for Clk_period;
Addr <= "1011000001110";
Trees_din <= "00000011000000000011011000000100";
wait for Clk_period;
Addr <= "1011000001111";
Trees_din <= "00000000010110010101100001000101";
wait for Clk_period;
Addr <= "1011000010000";
Trees_din <= "00000000001100110101100001000101";
wait for Clk_period;



----------tree 44-------------------

Addr <= "1011000010001";
Trees_din <= "00000101000000000010111110000000";
wait for Clk_period;
Addr <= "1011000010010";
Trees_din <= "00000110000000000100000001000000";
wait for Clk_period;
Addr <= "1011000010011";
Trees_din <= "00000101000000000010000100100000";
wait for Clk_period;
Addr <= "1011000010100";
Trees_din <= "00000111000000000100011000010000";
wait for Clk_period;
Addr <= "1011000010101";
Trees_din <= "00000000000000000001101100001000";
wait for Clk_period;
Addr <= "1011000010110";
Trees_din <= "00000111000000000011100100000100";
wait for Clk_period;
Addr <= "1011000010111";
Trees_din <= "00000000001000000000000000000011";
wait for Clk_period;
Addr <= "1011000011000";
Trees_din <= "00000000001000000000000000000011";
wait for Clk_period;
Addr <= "1011000011001";
Trees_din <= "00000100000000000011101100000100";
wait for Clk_period;
Addr <= "1011000011010";
Trees_din <= "00000000011000000000000000000011";
wait for Clk_period;
Addr <= "1011000011011";
Trees_din <= "00000000000010010000000000000011";
wait for Clk_period;
Addr <= "1011000011100";
Trees_din <= "00000000000000000110000000001000";
wait for Clk_period;
Addr <= "1011000011101";
Trees_din <= "00000001000000000010110000000100";
wait for Clk_period;
Addr <= "1011000011110";
Trees_din <= "00000000001101100000000000000011";
wait for Clk_period;
Addr <= "1011000011111";
Trees_din <= "00000000010101100000000000000011";
wait for Clk_period;
Addr <= "1011000100000";
Trees_din <= "00000100000000000001001000000100";
wait for Clk_period;
Addr <= "1011000100001";
Trees_din <= "00000000010000100000000000000011";
wait for Clk_period;
Addr <= "1011000100010";
Trees_din <= "00000000010010010000000000000011";
wait for Clk_period;
Addr <= "1011000100011";
Trees_din <= "00000110000000000011001100010000";
wait for Clk_period;
Addr <= "1011000100100";
Trees_din <= "00000111000000000000101000001000";
wait for Clk_period;
Addr <= "1011000100101";
Trees_din <= "00000010000000000010010000000100";
wait for Clk_period;
Addr <= "1011000100110";
Trees_din <= "00000000001100000000000000000011";
wait for Clk_period;
Addr <= "1011000100111";
Trees_din <= "00000000001101000000000000000011";
wait for Clk_period;
Addr <= "1011000101000";
Trees_din <= "00000010000000000011010000000100";
wait for Clk_period;
Addr <= "1011000101001";
Trees_din <= "00000000000010110000000000000011";
wait for Clk_period;
Addr <= "1011000101010";
Trees_din <= "00000000001110010000000000000011";
wait for Clk_period;
Addr <= "1011000101011";
Trees_din <= "00000000000000000000001100001000";
wait for Clk_period;
Addr <= "1011000101100";
Trees_din <= "00000110000000000011001100000100";
wait for Clk_period;
Addr <= "1011000101101";
Trees_din <= "00000000010010110000000000000011";
wait for Clk_period;
Addr <= "1011000101110";
Trees_din <= "00000000001100000000000000000011";
wait for Clk_period;
Addr <= "1011000101111";
Trees_din <= "00000101000000000101010000000100";
wait for Clk_period;
Addr <= "1011000110000";
Trees_din <= "00000000010110010000000000000011";
wait for Clk_period;
Addr <= "1011000110001";
Trees_din <= "00000000001001000000000000000011";
wait for Clk_period;
Addr <= "1011000110010";
Trees_din <= "00000100000000000100000100100000";
wait for Clk_period;
Addr <= "1011000110011";
Trees_din <= "00000000000000000001010000010000";
wait for Clk_period;
Addr <= "1011000110100";
Trees_din <= "00000011000000000011111100001000";
wait for Clk_period;
Addr <= "1011000110101";
Trees_din <= "00000001000000000001110000000100";
wait for Clk_period;
Addr <= "1011000110110";
Trees_din <= "00000000000111110000000000000011";
wait for Clk_period;
Addr <= "1011000110111";
Trees_din <= "00000000010111110000000000000011";
wait for Clk_period;
Addr <= "1011000111000";
Trees_din <= "00000111000000000001011100000100";
wait for Clk_period;
Addr <= "1011000111001";
Trees_din <= "00000000000010000000000000000011";
wait for Clk_period;
Addr <= "1011000111010";
Trees_din <= "00000000011000000000000000000011";
wait for Clk_period;
Addr <= "1011000111011";
Trees_din <= "00000011000000000000110000001000";
wait for Clk_period;
Addr <= "1011000111100";
Trees_din <= "00000010000000000100010000000100";
wait for Clk_period;
Addr <= "1011000111101";
Trees_din <= "00000000001001010000000000000011";
wait for Clk_period;
Addr <= "1011000111110";
Trees_din <= "00000000000011100000000000000011";
wait for Clk_period;
Addr <= "1011000111111";
Trees_din <= "00000110000000000101101100000100";
wait for Clk_period;
Addr <= "1011001000000";
Trees_din <= "00000000010100010000000000000011";
wait for Clk_period;
Addr <= "1011001000001";
Trees_din <= "00000000011000100000000000000011";
wait for Clk_period;
Addr <= "1011001000010";
Trees_din <= "00000011000000000100111100010000";
wait for Clk_period;
Addr <= "1011001000011";
Trees_din <= "00000111000000000001010000001000";
wait for Clk_period;
Addr <= "1011001000100";
Trees_din <= "00000010000000000101101000000100";
wait for Clk_period;
Addr <= "1011001000101";
Trees_din <= "00000000010100010000000000000011";
wait for Clk_period;
Addr <= "1011001000110";
Trees_din <= "00000000001101000000000000000011";
wait for Clk_period;
Addr <= "1011001000111";
Trees_din <= "00000000000000000110010000000100";
wait for Clk_period;
Addr <= "1011001001000";
Trees_din <= "00000000000101100000000000000011";
wait for Clk_period;
Addr <= "1011001001001";
Trees_din <= "00000000010100000000000000000011";
wait for Clk_period;
Addr <= "1011001001010";
Trees_din <= "00000101000000000011111100001000";
wait for Clk_period;
Addr <= "1011001001011";
Trees_din <= "00000111000000000000111000000100";
wait for Clk_period;
Addr <= "1011001001100";
Trees_din <= "00000000000000000000000000000011";
wait for Clk_period;
Addr <= "1011001001101";
Trees_din <= "00000000000110110000000000000011";
wait for Clk_period;
Addr <= "1011001001110";
Trees_din <= "00000011000000000101000000000100";
wait for Clk_period;
Addr <= "1011001001111";
Trees_din <= "00000000001001100000000000000011";
wait for Clk_period;
Addr <= "1011001010000";
Trees_din <= "00000000010011100000000000000011";
wait for Clk_period;
Addr <= "1011001010001";
Trees_din <= "00000011000000000101000101000000";
wait for Clk_period;
Addr <= "1011001010010";
Trees_din <= "00000110000000000011101000100000";
wait for Clk_period;
Addr <= "1011001010011";
Trees_din <= "00000111000000000000001100010000";
wait for Clk_period;
Addr <= "1011001010100";
Trees_din <= "00000010000000000000011100001000";
wait for Clk_period;
Addr <= "1011001010101";
Trees_din <= "00000100000000000000100000000100";
wait for Clk_period;
Addr <= "1011001010110";
Trees_din <= "00000000010111000000000000000011";
wait for Clk_period;
Addr <= "1011001010111";
Trees_din <= "00000000000000000000000000000011";
wait for Clk_period;
Addr <= "1011001011000";
Trees_din <= "00000001000000000100010100000100";
wait for Clk_period;
Addr <= "1011001011001";
Trees_din <= "00000000000000110000000000000011";
wait for Clk_period;
Addr <= "1011001011010";
Trees_din <= "00000000000010010000000000000011";
wait for Clk_period;
Addr <= "1011001011011";
Trees_din <= "00000011000000000010010000001000";
wait for Clk_period;
Addr <= "1011001011100";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "1011001011101";
Trees_din <= "00000000001001000000000000000011";
wait for Clk_period;
Addr <= "1011001011110";
Trees_din <= "00000000001010110000000000000011";
wait for Clk_period;
Addr <= "1011001011111";
Trees_din <= "00000111000000000100101000000100";
wait for Clk_period;
Addr <= "1011001100000";
Trees_din <= "00000000010110110000000000000011";
wait for Clk_period;
Addr <= "1011001100001";
Trees_din <= "00000000001101110000000000000011";
wait for Clk_period;
Addr <= "1011001100010";
Trees_din <= "00000111000000000100000000010000";
wait for Clk_period;
Addr <= "1011001100011";
Trees_din <= "00000000000000000100001100001000";
wait for Clk_period;
Addr <= "1011001100100";
Trees_din <= "00000111000000000010100000000100";
wait for Clk_period;
Addr <= "1011001100101";
Trees_din <= "00000000000001000000000000000011";
wait for Clk_period;
Addr <= "1011001100110";
Trees_din <= "00000000001100010000000000000011";
wait for Clk_period;
Addr <= "1011001100111";
Trees_din <= "00000000000000000100001000000100";
wait for Clk_period;
Addr <= "1011001101000";
Trees_din <= "00000000001000000000000000000011";
wait for Clk_period;
Addr <= "1011001101001";
Trees_din <= "00000000010000100000000000000011";
wait for Clk_period;
Addr <= "1011001101010";
Trees_din <= "00000010000000000000010000001000";
wait for Clk_period;
Addr <= "1011001101011";
Trees_din <= "00000110000000000100100100000100";
wait for Clk_period;
Addr <= "1011001101100";
Trees_din <= "00000000010101010000000000000011";
wait for Clk_period;
Addr <= "1011001101101";
Trees_din <= "00000000010100110000000000000011";
wait for Clk_period;
Addr <= "1011001101110";
Trees_din <= "00000110000000000001111000000100";
wait for Clk_period;
Addr <= "1011001101111";
Trees_din <= "00000000001110000000000000000011";
wait for Clk_period;
Addr <= "1011001110000";
Trees_din <= "00000000001000010000000000000011";
wait for Clk_period;
Addr <= "1011001110001";
Trees_din <= "00000101000000000101100000100000";
wait for Clk_period;
Addr <= "1011001110010";
Trees_din <= "00000110000000000001110000010000";
wait for Clk_period;
Addr <= "1011001110011";
Trees_din <= "00000100000000000100100000001000";
wait for Clk_period;
Addr <= "1011001110100";
Trees_din <= "00000000000000000011011000000100";
wait for Clk_period;
Addr <= "1011001110101";
Trees_din <= "00000000001101010000000000000011";
wait for Clk_period;
Addr <= "1011001110110";
Trees_din <= "00000000001010000000000000000011";
wait for Clk_period;
Addr <= "1011001110111";
Trees_din <= "00000110000000000101111000000100";
wait for Clk_period;
Addr <= "1011001111000";
Trees_din <= "00000000001010100000000000000011";
wait for Clk_period;
Addr <= "1011001111001";
Trees_din <= "00000000010100100000000000000011";
wait for Clk_period;
Addr <= "1011001111010";
Trees_din <= "00000111000000000000010100001000";
wait for Clk_period;
Addr <= "1011001111011";
Trees_din <= "00000100000000000010110000000100";
wait for Clk_period;
Addr <= "1011001111100";
Trees_din <= "00000000010011010000000000000011";
wait for Clk_period;
Addr <= "1011001111101";
Trees_din <= "00000000001110100000000000000011";
wait for Clk_period;
Addr <= "1011001111110";
Trees_din <= "00000010000000000010110000000100";
wait for Clk_period;
Addr <= "1011001111111";
Trees_din <= "00000000001111010000000000000011";
wait for Clk_period;
Addr <= "1011010000000";
Trees_din <= "00000000000111010000000000000011";
wait for Clk_period;
Addr <= "1011010000001";
Trees_din <= "00000000000000000000111100010000";
wait for Clk_period;
Addr <= "1011010000010";
Trees_din <= "00000001000000000010000000001000";
wait for Clk_period;
Addr <= "1011010000011";
Trees_din <= "00000000000000000101110000000100";
wait for Clk_period;
Addr <= "1011010000100";
Trees_din <= "00000000010000100000000000000011";
wait for Clk_period;
Addr <= "1011010000101";
Trees_din <= "00000000000011110000000000000011";
wait for Clk_period;
Addr <= "1011010000110";
Trees_din <= "00000011000000000001111000000100";
wait for Clk_period;
Addr <= "1011010000111";
Trees_din <= "00000000001011110000000000000011";
wait for Clk_period;
Addr <= "1011010001000";
Trees_din <= "00000000010110010000000000000011";
wait for Clk_period;
Addr <= "1011010001001";
Trees_din <= "00000010000000000100010100001000";
wait for Clk_period;
Addr <= "1011010001010";
Trees_din <= "00000110000000000001111000000100";
wait for Clk_period;
Addr <= "1011010001011";
Trees_din <= "00000000000001100000000000000011";
wait for Clk_period;
Addr <= "1011010001100";
Trees_din <= "00000000000000110000000000000011";
wait for Clk_period;
Addr <= "1011010001101";
Trees_din <= "00000100000000000100001000000100";
wait for Clk_period;
Addr <= "1011010001110";
Trees_din <= "00000000010001100000000000000011";
wait for Clk_period;
Addr <= "1011010001111";
Trees_din <= "00000000010110000000000000000011";
wait for Clk_period;



----------tree 45-------------------

Addr <= "1011010010000";
Trees_din <= "00000111000000000101000110000000";
wait for Clk_period;
Addr <= "1011010010001";
Trees_din <= "00000101000000000010111101000000";
wait for Clk_period;
Addr <= "1011010010010";
Trees_din <= "00000110000000000011100100100000";
wait for Clk_period;
Addr <= "1011010010011";
Trees_din <= "00000100000000000001100100010000";
wait for Clk_period;
Addr <= "1011010010100";
Trees_din <= "00000011000000000101111100001000";
wait for Clk_period;
Addr <= "1011010010101";
Trees_din <= "00000110000000000001011000000100";
wait for Clk_period;
Addr <= "1011010010110";
Trees_din <= "00000000000111110101110000111101";
wait for Clk_period;
Addr <= "1011010010111";
Trees_din <= "00000000010101000101110000111101";
wait for Clk_period;
Addr <= "1011010011000";
Trees_din <= "00000001000000000100101000000100";
wait for Clk_period;
Addr <= "1011010011001";
Trees_din <= "00000000000101110101110000111101";
wait for Clk_period;
Addr <= "1011010011010";
Trees_din <= "00000000010110010101110000111101";
wait for Clk_period;
Addr <= "1011010011011";
Trees_din <= "00000011000000000010010000001000";
wait for Clk_period;
Addr <= "1011010011100";
Trees_din <= "00000110000000000000111100000100";
wait for Clk_period;
Addr <= "1011010011101";
Trees_din <= "00000000010111100101110000111101";
wait for Clk_period;
Addr <= "1011010011110";
Trees_din <= "00000000010100100101110000111101";
wait for Clk_period;
Addr <= "1011010011111";
Trees_din <= "00000010000000000101000100000100";
wait for Clk_period;
Addr <= "1011010100000";
Trees_din <= "00000000000101000101110000111101";
wait for Clk_period;
Addr <= "1011010100001";
Trees_din <= "00000000000011000101110000111101";
wait for Clk_period;
Addr <= "1011010100010";
Trees_din <= "00000100000000000010010100010000";
wait for Clk_period;
Addr <= "1011010100011";
Trees_din <= "00000110000000000011101000001000";
wait for Clk_period;
Addr <= "1011010100100";
Trees_din <= "00000110000000000010001000000100";
wait for Clk_period;
Addr <= "1011010100101";
Trees_din <= "00000000001011000101110000111101";
wait for Clk_period;
Addr <= "1011010100110";
Trees_din <= "00000000000111100101110000111101";
wait for Clk_period;
Addr <= "1011010100111";
Trees_din <= "00000011000000000101010000000100";
wait for Clk_period;
Addr <= "1011010101000";
Trees_din <= "00000000000101000101110000111101";
wait for Clk_period;
Addr <= "1011010101001";
Trees_din <= "00000000001100110101110000111101";
wait for Clk_period;
Addr <= "1011010101010";
Trees_din <= "00000010000000000001001000001000";
wait for Clk_period;
Addr <= "1011010101011";
Trees_din <= "00000001000000000011101100000100";
wait for Clk_period;
Addr <= "1011010101100";
Trees_din <= "00000000000101010101110000111101";
wait for Clk_period;
Addr <= "1011010101101";
Trees_din <= "00000000000001100101110000111101";
wait for Clk_period;
Addr <= "1011010101110";
Trees_din <= "00000110000000000101001100000100";
wait for Clk_period;
Addr <= "1011010101111";
Trees_din <= "00000000001010000101110000111101";
wait for Clk_period;
Addr <= "1011010110000";
Trees_din <= "00000000010011100101110000111101";
wait for Clk_period;
Addr <= "1011010110001";
Trees_din <= "00000110000000000010111100100000";
wait for Clk_period;
Addr <= "1011010110010";
Trees_din <= "00000001000000000101111100010000";
wait for Clk_period;
Addr <= "1011010110011";
Trees_din <= "00000010000000000000100000001000";
wait for Clk_period;
Addr <= "1011010110100";
Trees_din <= "00000011000000000000011000000100";
wait for Clk_period;
Addr <= "1011010110101";
Trees_din <= "00000000001011000101110000111101";
wait for Clk_period;
Addr <= "1011010110110";
Trees_din <= "00000000001000010101110000111101";
wait for Clk_period;
Addr <= "1011010110111";
Trees_din <= "00000011000000000110000000000100";
wait for Clk_period;
Addr <= "1011010111000";
Trees_din <= "00000000000000010101110000111101";
wait for Clk_period;
Addr <= "1011010111001";
Trees_din <= "00000000001100110101110000111101";
wait for Clk_period;
Addr <= "1011010111010";
Trees_din <= "00000101000000000011111100001000";
wait for Clk_period;
Addr <= "1011010111011";
Trees_din <= "00000100000000000000010000000100";
wait for Clk_period;
Addr <= "1011010111100";
Trees_din <= "00000000001111000101110000111101";
wait for Clk_period;
Addr <= "1011010111101";
Trees_din <= "00000000001000000101110000111101";
wait for Clk_period;
Addr <= "1011010111110";
Trees_din <= "00000111000000000101101100000100";
wait for Clk_period;
Addr <= "1011010111111";
Trees_din <= "00000000000101010101110000111101";
wait for Clk_period;
Addr <= "1011011000000";
Trees_din <= "00000000000011100101110000111101";
wait for Clk_period;
Addr <= "1011011000001";
Trees_din <= "00000100000000000011110000010000";
wait for Clk_period;
Addr <= "1011011000010";
Trees_din <= "00000000000000000100000100001000";
wait for Clk_period;
Addr <= "1011011000011";
Trees_din <= "00000110000000000000011100000100";
wait for Clk_period;
Addr <= "1011011000100";
Trees_din <= "00000000001011110101110000111101";
wait for Clk_period;
Addr <= "1011011000101";
Trees_din <= "00000000000001110101110000111101";
wait for Clk_period;
Addr <= "1011011000110";
Trees_din <= "00000110000000000110010000000100";
wait for Clk_period;
Addr <= "1011011000111";
Trees_din <= "00000000001010000101110000111101";
wait for Clk_period;
Addr <= "1011011001000";
Trees_din <= "00000000000010010101110000111101";
wait for Clk_period;
Addr <= "1011011001001";
Trees_din <= "00000111000000000100001100001000";
wait for Clk_period;
Addr <= "1011011001010";
Trees_din <= "00000000000000000001110100000100";
wait for Clk_period;
Addr <= "1011011001011";
Trees_din <= "00000000010011010101110000111101";
wait for Clk_period;
Addr <= "1011011001100";
Trees_din <= "00000000010110110101110000111101";
wait for Clk_period;
Addr <= "1011011001101";
Trees_din <= "00000001000000000000110100000100";
wait for Clk_period;
Addr <= "1011011001110";
Trees_din <= "00000000001100000101110000111101";
wait for Clk_period;
Addr <= "1011011001111";
Trees_din <= "00000000000001000101110000111101";
wait for Clk_period;
Addr <= "1011011010000";
Trees_din <= "00000110000000000101100001000000";
wait for Clk_period;
Addr <= "1011011010001";
Trees_din <= "00000111000000000001101000100000";
wait for Clk_period;
Addr <= "1011011010010";
Trees_din <= "00000001000000000000011100010000";
wait for Clk_period;
Addr <= "1011011010011";
Trees_din <= "00000110000000000110001100001000";
wait for Clk_period;
Addr <= "1011011010100";
Trees_din <= "00000111000000000101001100000100";
wait for Clk_period;
Addr <= "1011011010101";
Trees_din <= "00000000010110000101110000111101";
wait for Clk_period;
Addr <= "1011011010110";
Trees_din <= "00000000010101010101110000111101";
wait for Clk_period;
Addr <= "1011011010111";
Trees_din <= "00000010000000000101010000000100";
wait for Clk_period;
Addr <= "1011011011000";
Trees_din <= "00000000001001000101110000111101";
wait for Clk_period;
Addr <= "1011011011001";
Trees_din <= "00000000010111010101110000111101";
wait for Clk_period;
Addr <= "1011011011010";
Trees_din <= "00000000000000000101100000001000";
wait for Clk_period;
Addr <= "1011011011011";
Trees_din <= "00000111000000000011110100000100";
wait for Clk_period;
Addr <= "1011011011100";
Trees_din <= "00000000010100100101110000111101";
wait for Clk_period;
Addr <= "1011011011101";
Trees_din <= "00000000000001010101110000111101";
wait for Clk_period;
Addr <= "1011011011110";
Trees_din <= "00000110000000000100001000000100";
wait for Clk_period;
Addr <= "1011011011111";
Trees_din <= "00000000010101000101110000111101";
wait for Clk_period;
Addr <= "1011011100000";
Trees_din <= "00000000001011000101110000111101";
wait for Clk_period;
Addr <= "1011011100001";
Trees_din <= "00000011000000000100001100010000";
wait for Clk_period;
Addr <= "1011011100010";
Trees_din <= "00000000000000000001110100001000";
wait for Clk_period;
Addr <= "1011011100011";
Trees_din <= "00000110000000000001011000000100";
wait for Clk_period;
Addr <= "1011011100100";
Trees_din <= "00000000000011100101110000111101";
wait for Clk_period;
Addr <= "1011011100101";
Trees_din <= "00000000001011010101110000111101";
wait for Clk_period;
Addr <= "1011011100110";
Trees_din <= "00000110000000000001000100000100";
wait for Clk_period;
Addr <= "1011011100111";
Trees_din <= "00000000000010010101110000111101";
wait for Clk_period;
Addr <= "1011011101000";
Trees_din <= "00000000001101110101110000111101";
wait for Clk_period;
Addr <= "1011011101001";
Trees_din <= "00000100000000000000001000001000";
wait for Clk_period;
Addr <= "1011011101010";
Trees_din <= "00000010000000000101011000000100";
wait for Clk_period;
Addr <= "1011011101011";
Trees_din <= "00000000001100100101110000111101";
wait for Clk_period;
Addr <= "1011011101100";
Trees_din <= "00000000001111000101110000111101";
wait for Clk_period;
Addr <= "1011011101101";
Trees_din <= "00000101000000000001011000000100";
wait for Clk_period;
Addr <= "1011011101110";
Trees_din <= "00000000000010010101110000111101";
wait for Clk_period;
Addr <= "1011011101111";
Trees_din <= "00000000000111100101110000111101";
wait for Clk_period;
Addr <= "1011011110000";
Trees_din <= "00000110000000000101001100100000";
wait for Clk_period;
Addr <= "1011011110001";
Trees_din <= "00000101000000000100100100010000";
wait for Clk_period;
Addr <= "1011011110010";
Trees_din <= "00000110000000000100100000001000";
wait for Clk_period;
Addr <= "1011011110011";
Trees_din <= "00000110000000000001010100000100";
wait for Clk_period;
Addr <= "1011011110100";
Trees_din <= "00000000010111010101110000111101";
wait for Clk_period;
Addr <= "1011011110101";
Trees_din <= "00000000010010100101110000111101";
wait for Clk_period;
Addr <= "1011011110110";
Trees_din <= "00000011000000000100110000000100";
wait for Clk_period;
Addr <= "1011011110111";
Trees_din <= "00000000000101100101110000111101";
wait for Clk_period;
Addr <= "1011011111000";
Trees_din <= "00000000001111000101110000111101";
wait for Clk_period;
Addr <= "1011011111001";
Trees_din <= "00000001000000000001000100001000";
wait for Clk_period;
Addr <= "1011011111010";
Trees_din <= "00000110000000000101101000000100";
wait for Clk_period;
Addr <= "1011011111011";
Trees_din <= "00000000010111000101110000111101";
wait for Clk_period;
Addr <= "1011011111100";
Trees_din <= "00000000000100110101110000111101";
wait for Clk_period;
Addr <= "1011011111101";
Trees_din <= "00000000000000000000110100000100";
wait for Clk_period;
Addr <= "1011011111110";
Trees_din <= "00000000001111010101110000111101";
wait for Clk_period;
Addr <= "1011011111111";
Trees_din <= "00000000000110110101110000111101";
wait for Clk_period;
Addr <= "1011100000000";
Trees_din <= "00000101000000000100000000010000";
wait for Clk_period;
Addr <= "1011100000001";
Trees_din <= "00000000000000000010100000001000";
wait for Clk_period;
Addr <= "1011100000010";
Trees_din <= "00000100000000000101100000000100";
wait for Clk_period;
Addr <= "1011100000011";
Trees_din <= "00000000011001000101110000111101";
wait for Clk_period;
Addr <= "1011100000100";
Trees_din <= "00000000001001010101110000111101";
wait for Clk_period;
Addr <= "1011100000101";
Trees_din <= "00000111000000000010010000000100";
wait for Clk_period;
Addr <= "1011100000110";
Trees_din <= "00000000001010110101110000111101";
wait for Clk_period;
Addr <= "1011100000111";
Trees_din <= "00000000000011110101110000111101";
wait for Clk_period;
Addr <= "1011100001000";
Trees_din <= "00000110000000000011001100001000";
wait for Clk_period;
Addr <= "1011100001001";
Trees_din <= "00000111000000000000010100000100";
wait for Clk_period;
Addr <= "1011100001010";
Trees_din <= "00000000011000000101110000111101";
wait for Clk_period;
Addr <= "1011100001011";
Trees_din <= "00000000001010100101110000111101";
wait for Clk_period;
Addr <= "1011100001100";
Trees_din <= "00000100000000000000011000000100";
wait for Clk_period;
Addr <= "1011100001101";
Trees_din <= "00000000010111000101110000111101";
wait for Clk_period;
Addr <= "1011100001110";
Trees_din <= "00000000000000010101110000111101";
wait for Clk_period;



----------tree 46-------------------

Addr <= "1011100001111";
Trees_din <= "00000010000000000101000110000000";
wait for Clk_period;
Addr <= "1011100010000";
Trees_din <= "00000001000000000101110001000000";
wait for Clk_period;
Addr <= "1011100010001";
Trees_din <= "00000110000000000001111100100000";
wait for Clk_period;
Addr <= "1011100010010";
Trees_din <= "00000111000000000000101100010000";
wait for Clk_period;
Addr <= "1011100010011";
Trees_din <= "00000010000000000011001000001000";
wait for Clk_period;
Addr <= "1011100010100";
Trees_din <= "00000000000000000001101100000100";
wait for Clk_period;
Addr <= "1011100010101";
Trees_din <= "00000000010000110101111000111001";
wait for Clk_period;
Addr <= "1011100010110";
Trees_din <= "00000000001010010101111000111001";
wait for Clk_period;
Addr <= "1011100010111";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "1011100011000";
Trees_din <= "00000000000100010101111000111001";
wait for Clk_period;
Addr <= "1011100011001";
Trees_din <= "00000000010101110101111000111001";
wait for Clk_period;
Addr <= "1011100011010";
Trees_din <= "00000101000000000000001100001000";
wait for Clk_period;
Addr <= "1011100011011";
Trees_din <= "00000000000000000001010000000100";
wait for Clk_period;
Addr <= "1011100011100";
Trees_din <= "00000000001101010101111000111001";
wait for Clk_period;
Addr <= "1011100011101";
Trees_din <= "00000000001111000101111000111001";
wait for Clk_period;
Addr <= "1011100011110";
Trees_din <= "00000010000000000001101100000100";
wait for Clk_period;
Addr <= "1011100011111";
Trees_din <= "00000000010000000101111000111001";
wait for Clk_period;
Addr <= "1011100100000";
Trees_din <= "00000000010110110101111000111001";
wait for Clk_period;
Addr <= "1011100100001";
Trees_din <= "00000100000000000011011100010000";
wait for Clk_period;
Addr <= "1011100100010";
Trees_din <= "00000000000000000000000000001000";
wait for Clk_period;
Addr <= "1011100100011";
Trees_din <= "00000011000000000011111100000100";
wait for Clk_period;
Addr <= "1011100100100";
Trees_din <= "00000000000000100101111000111001";
wait for Clk_period;
Addr <= "1011100100101";
Trees_din <= "00000000000001110101111000111001";
wait for Clk_period;
Addr <= "1011100100110";
Trees_din <= "00000000000000000101001000000100";
wait for Clk_period;
Addr <= "1011100100111";
Trees_din <= "00000000010010110101111000111001";
wait for Clk_period;
Addr <= "1011100101000";
Trees_din <= "00000000010110110101111000111001";
wait for Clk_period;
Addr <= "1011100101001";
Trees_din <= "00000101000000000010000000001000";
wait for Clk_period;
Addr <= "1011100101010";
Trees_din <= "00000001000000000100010100000100";
wait for Clk_period;
Addr <= "1011100101011";
Trees_din <= "00000000010010100101111000111001";
wait for Clk_period;
Addr <= "1011100101100";
Trees_din <= "00000000010101000101111000111001";
wait for Clk_period;
Addr <= "1011100101101";
Trees_din <= "00000001000000000110001100000100";
wait for Clk_period;
Addr <= "1011100101110";
Trees_din <= "00000000000011010101111000111001";
wait for Clk_period;
Addr <= "1011100101111";
Trees_din <= "00000000000100010101111000111001";
wait for Clk_period;
Addr <= "1011100110000";
Trees_din <= "00000101000000000100101100100000";
wait for Clk_period;
Addr <= "1011100110001";
Trees_din <= "00000001000000000100011100010000";
wait for Clk_period;
Addr <= "1011100110010";
Trees_din <= "00000000000000000010010100001000";
wait for Clk_period;
Addr <= "1011100110011";
Trees_din <= "00000101000000000101001000000100";
wait for Clk_period;
Addr <= "1011100110100";
Trees_din <= "00000000001011110101111000111001";
wait for Clk_period;
Addr <= "1011100110101";
Trees_din <= "00000000001100000101111000111001";
wait for Clk_period;
Addr <= "1011100110110";
Trees_din <= "00000011000000000101011100000100";
wait for Clk_period;
Addr <= "1011100110111";
Trees_din <= "00000000001001010101111000111001";
wait for Clk_period;
Addr <= "1011100111000";
Trees_din <= "00000000000011010101111000111001";
wait for Clk_period;
Addr <= "1011100111001";
Trees_din <= "00000001000000000100001100001000";
wait for Clk_period;
Addr <= "1011100111010";
Trees_din <= "00000010000000000010001100000100";
wait for Clk_period;
Addr <= "1011100111011";
Trees_din <= "00000000001111100101111000111001";
wait for Clk_period;
Addr <= "1011100111100";
Trees_din <= "00000000000100110101111000111001";
wait for Clk_period;
Addr <= "1011100111101";
Trees_din <= "00000000000000000101001100000100";
wait for Clk_period;
Addr <= "1011100111110";
Trees_din <= "00000000001001100101111000111001";
wait for Clk_period;
Addr <= "1011100111111";
Trees_din <= "00000000010101100101111000111001";
wait for Clk_period;
Addr <= "1011101000000";
Trees_din <= "00000110000000000001010100010000";
wait for Clk_period;
Addr <= "1011101000001";
Trees_din <= "00000010000000000000011100001000";
wait for Clk_period;
Addr <= "1011101000010";
Trees_din <= "00000001000000000001001100000100";
wait for Clk_period;
Addr <= "1011101000011";
Trees_din <= "00000000010111110101111000111001";
wait for Clk_period;
Addr <= "1011101000100";
Trees_din <= "00000000010010000101111000111001";
wait for Clk_period;
Addr <= "1011101000101";
Trees_din <= "00000101000000000010111000000100";
wait for Clk_period;
Addr <= "1011101000110";
Trees_din <= "00000000000010000101111000111001";
wait for Clk_period;
Addr <= "1011101000111";
Trees_din <= "00000000010101000101111000111001";
wait for Clk_period;
Addr <= "1011101001000";
Trees_din <= "00000010000000000000011000001000";
wait for Clk_period;
Addr <= "1011101001001";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "1011101001010";
Trees_din <= "00000000000011110101111000111001";
wait for Clk_period;
Addr <= "1011101001011";
Trees_din <= "00000000010110110101111000111001";
wait for Clk_period;
Addr <= "1011101001100";
Trees_din <= "00000110000000000011110100000100";
wait for Clk_period;
Addr <= "1011101001101";
Trees_din <= "00000000010010100101111000111001";
wait for Clk_period;
Addr <= "1011101001110";
Trees_din <= "00000000001010110101111000111001";
wait for Clk_period;
Addr <= "1011101001111";
Trees_din <= "00000011000000000011100001000000";
wait for Clk_period;
Addr <= "1011101010000";
Trees_din <= "00000100000000000011110100100000";
wait for Clk_period;
Addr <= "1011101010001";
Trees_din <= "00000010000000000101011000010000";
wait for Clk_period;
Addr <= "1011101010010";
Trees_din <= "00000000000000000010010100001000";
wait for Clk_period;
Addr <= "1011101010011";
Trees_din <= "00000000000000000010111100000100";
wait for Clk_period;
Addr <= "1011101010100";
Trees_din <= "00000000010011000101111000111001";
wait for Clk_period;
Addr <= "1011101010101";
Trees_din <= "00000000000111110101111000111001";
wait for Clk_period;
Addr <= "1011101010110";
Trees_din <= "00000100000000000001010000000100";
wait for Clk_period;
Addr <= "1011101010111";
Trees_din <= "00000000010010110101111000111001";
wait for Clk_period;
Addr <= "1011101011000";
Trees_din <= "00000000001001000101111000111001";
wait for Clk_period;
Addr <= "1011101011001";
Trees_din <= "00000101000000000001101100001000";
wait for Clk_period;
Addr <= "1011101011010";
Trees_din <= "00000111000000000001110100000100";
wait for Clk_period;
Addr <= "1011101011011";
Trees_din <= "00000000010111000101111000111001";
wait for Clk_period;
Addr <= "1011101011100";
Trees_din <= "00000000001000110101111000111001";
wait for Clk_period;
Addr <= "1011101011101";
Trees_din <= "00000000000000000101100100000100";
wait for Clk_period;
Addr <= "1011101011110";
Trees_din <= "00000000001101010101111000111001";
wait for Clk_period;
Addr <= "1011101011111";
Trees_din <= "00000000001001100101111000111001";
wait for Clk_period;
Addr <= "1011101100000";
Trees_din <= "00000010000000000000001100010000";
wait for Clk_period;
Addr <= "1011101100001";
Trees_din <= "00000100000000000100111100001000";
wait for Clk_period;
Addr <= "1011101100010";
Trees_din <= "00000010000000000010111000000100";
wait for Clk_period;
Addr <= "1011101100011";
Trees_din <= "00000000010011100101111000111001";
wait for Clk_period;
Addr <= "1011101100100";
Trees_din <= "00000000001010100101111000111001";
wait for Clk_period;
Addr <= "1011101100101";
Trees_din <= "00000101000000000110001000000100";
wait for Clk_period;
Addr <= "1011101100110";
Trees_din <= "00000000000011000101111000111001";
wait for Clk_period;
Addr <= "1011101100111";
Trees_din <= "00000000001000110101111000111001";
wait for Clk_period;
Addr <= "1011101101000";
Trees_din <= "00000111000000000100010100001000";
wait for Clk_period;
Addr <= "1011101101001";
Trees_din <= "00000001000000000101100100000100";
wait for Clk_period;
Addr <= "1011101101010";
Trees_din <= "00000000000010000101111000111001";
wait for Clk_period;
Addr <= "1011101101011";
Trees_din <= "00000000000101000101111000111001";
wait for Clk_period;
Addr <= "1011101101100";
Trees_din <= "00000001000000000001111100000100";
wait for Clk_period;
Addr <= "1011101101101";
Trees_din <= "00000000010000110101111000111001";
wait for Clk_period;
Addr <= "1011101101110";
Trees_din <= "00000000000001000101111000111001";
wait for Clk_period;
Addr <= "1011101101111";
Trees_din <= "00000100000000000100001000100000";
wait for Clk_period;
Addr <= "1011101110000";
Trees_din <= "00000001000000000001101000010000";
wait for Clk_period;
Addr <= "1011101110001";
Trees_din <= "00000111000000000000111000001000";
wait for Clk_period;
Addr <= "1011101110010";
Trees_din <= "00000101000000000100101000000100";
wait for Clk_period;
Addr <= "1011101110011";
Trees_din <= "00000000000011100101111000111001";
wait for Clk_period;
Addr <= "1011101110100";
Trees_din <= "00000000000000010101111000111001";
wait for Clk_period;
Addr <= "1011101110101";
Trees_din <= "00000001000000000001101000000100";
wait for Clk_period;
Addr <= "1011101110110";
Trees_din <= "00000000010000110101111000111001";
wait for Clk_period;
Addr <= "1011101110111";
Trees_din <= "00000000001101110101111000111001";
wait for Clk_period;
Addr <= "1011101111000";
Trees_din <= "00000000000000000001100000001000";
wait for Clk_period;
Addr <= "1011101111001";
Trees_din <= "00000110000000000001000000000100";
wait for Clk_period;
Addr <= "1011101111010";
Trees_din <= "00000000001011000101111000111001";
wait for Clk_period;
Addr <= "1011101111011";
Trees_din <= "00000000001101100101111000111001";
wait for Clk_period;
Addr <= "1011101111100";
Trees_din <= "00000100000000000100111000000100";
wait for Clk_period;
Addr <= "1011101111101";
Trees_din <= "00000000010101010101111000111001";
wait for Clk_period;
Addr <= "1011101111110";
Trees_din <= "00000000000000100101111000111001";
wait for Clk_period;
Addr <= "1011101111111";
Trees_din <= "00000010000000000000011000010000";
wait for Clk_period;
Addr <= "1011110000000";
Trees_din <= "00000010000000000100001000001000";
wait for Clk_period;
Addr <= "1011110000001";
Trees_din <= "00000001000000000100000100000100";
wait for Clk_period;
Addr <= "1011110000010";
Trees_din <= "00000000010100010101111000111001";
wait for Clk_period;
Addr <= "1011110000011";
Trees_din <= "00000000000100000101111000111001";
wait for Clk_period;
Addr <= "1011110000100";
Trees_din <= "00000011000000000101010000000100";
wait for Clk_period;
Addr <= "1011110000101";
Trees_din <= "00000000000010000101111000111001";
wait for Clk_period;
Addr <= "1011110000110";
Trees_din <= "00000000000111110101111000111001";
wait for Clk_period;
Addr <= "1011110000111";
Trees_din <= "00000111000000000011011100001000";
wait for Clk_period;
Addr <= "1011110001000";
Trees_din <= "00000000000000000001111000000100";
wait for Clk_period;
Addr <= "1011110001001";
Trees_din <= "00000000000000110101111000111001";
wait for Clk_period;
Addr <= "1011110001010";
Trees_din <= "00000000001001000101111000111001";
wait for Clk_period;
Addr <= "1011110001011";
Trees_din <= "00000011000000000010000000000100";
wait for Clk_period;
Addr <= "1011110001100";
Trees_din <= "00000000010110000101111000111001";
wait for Clk_period;
Addr <= "1011110001101";
Trees_din <= "00000000001100000101111000111001";
wait for Clk_period;



----------tree 47-------------------

Addr <= "1011110001110";
Trees_din <= "00000001000000000001000010000000";
wait for Clk_period;
Addr <= "1011110001111";
Trees_din <= "00000010000000000011100001000000";
wait for Clk_period;
Addr <= "1011110010000";
Trees_din <= "00000110000000000001001100100000";
wait for Clk_period;
Addr <= "1011110010001";
Trees_din <= "00000100000000000001110100010000";
wait for Clk_period;
Addr <= "1011110010010";
Trees_din <= "00000011000000000001010100001000";
wait for Clk_period;
Addr <= "1011110010011";
Trees_din <= "00000011000000000011110000000100";
wait for Clk_period;
Addr <= "1011110010100";
Trees_din <= "00000000010110100110000000110101";
wait for Clk_period;
Addr <= "1011110010101";
Trees_din <= "00000000001001000110000000110101";
wait for Clk_period;
Addr <= "1011110010110";
Trees_din <= "00000011000000000010011100000100";
wait for Clk_period;
Addr <= "1011110010111";
Trees_din <= "00000000001111110110000000110101";
wait for Clk_period;
Addr <= "1011110011000";
Trees_din <= "00000000001010100110000000110101";
wait for Clk_period;
Addr <= "1011110011001";
Trees_din <= "00000110000000000100111000001000";
wait for Clk_period;
Addr <= "1011110011010";
Trees_din <= "00000000000000000000110000000100";
wait for Clk_period;
Addr <= "1011110011011";
Trees_din <= "00000000001101010110000000110101";
wait for Clk_period;
Addr <= "1011110011100";
Trees_din <= "00000000010101110110000000110101";
wait for Clk_period;
Addr <= "1011110011101";
Trees_din <= "00000100000000000010011000000100";
wait for Clk_period;
Addr <= "1011110011110";
Trees_din <= "00000000010101000110000000110101";
wait for Clk_period;
Addr <= "1011110011111";
Trees_din <= "00000000010001010110000000110101";
wait for Clk_period;
Addr <= "1011110100000";
Trees_din <= "00000000000000000011110100010000";
wait for Clk_period;
Addr <= "1011110100001";
Trees_din <= "00000100000000000100010100001000";
wait for Clk_period;
Addr <= "1011110100010";
Trees_din <= "00000100000000000100100100000100";
wait for Clk_period;
Addr <= "1011110100011";
Trees_din <= "00000000001011100110000000110101";
wait for Clk_period;
Addr <= "1011110100100";
Trees_din <= "00000000000110010110000000110101";
wait for Clk_period;
Addr <= "1011110100101";
Trees_din <= "00000001000000000011111100000100";
wait for Clk_period;
Addr <= "1011110100110";
Trees_din <= "00000000001111100110000000110101";
wait for Clk_period;
Addr <= "1011110100111";
Trees_din <= "00000000010000100110000000110101";
wait for Clk_period;
Addr <= "1011110101000";
Trees_din <= "00000011000000000101101000001000";
wait for Clk_period;
Addr <= "1011110101001";
Trees_din <= "00000000000000000001111100000100";
wait for Clk_period;
Addr <= "1011110101010";
Trees_din <= "00000000011000000110000000110101";
wait for Clk_period;
Addr <= "1011110101011";
Trees_din <= "00000000000111100110000000110101";
wait for Clk_period;
Addr <= "1011110101100";
Trees_din <= "00000000000000000110001000000100";
wait for Clk_period;
Addr <= "1011110101101";
Trees_din <= "00000000001101000110000000110101";
wait for Clk_period;
Addr <= "1011110101110";
Trees_din <= "00000000000110110110000000110101";
wait for Clk_period;
Addr <= "1011110101111";
Trees_din <= "00000100000000000010110000100000";
wait for Clk_period;
Addr <= "1011110110000";
Trees_din <= "00000111000000000010101100010000";
wait for Clk_period;
Addr <= "1011110110001";
Trees_din <= "00000101000000000100011000001000";
wait for Clk_period;
Addr <= "1011110110010";
Trees_din <= "00000101000000000000001100000100";
wait for Clk_period;
Addr <= "1011110110011";
Trees_din <= "00000000000101100110000000110101";
wait for Clk_period;
Addr <= "1011110110100";
Trees_din <= "00000000000000110110000000110101";
wait for Clk_period;
Addr <= "1011110110101";
Trees_din <= "00000101000000000000110100000100";
wait for Clk_period;
Addr <= "1011110110110";
Trees_din <= "00000000001100100110000000110101";
wait for Clk_period;
Addr <= "1011110110111";
Trees_din <= "00000000001101010110000000110101";
wait for Clk_period;
Addr <= "1011110111000";
Trees_din <= "00000000000000000011101000001000";
wait for Clk_period;
Addr <= "1011110111001";
Trees_din <= "00000100000000000100110000000100";
wait for Clk_period;
Addr <= "1011110111010";
Trees_din <= "00000000010000100110000000110101";
wait for Clk_period;
Addr <= "1011110111011";
Trees_din <= "00000000010101010110000000110101";
wait for Clk_period;
Addr <= "1011110111100";
Trees_din <= "00000111000000000000101100000100";
wait for Clk_period;
Addr <= "1011110111101";
Trees_din <= "00000000010000110110000000110101";
wait for Clk_period;
Addr <= "1011110111110";
Trees_din <= "00000000010001110110000000110101";
wait for Clk_period;
Addr <= "1011110111111";
Trees_din <= "00000101000000000000001100010000";
wait for Clk_period;
Addr <= "1011111000000";
Trees_din <= "00000000000000000011111100001000";
wait for Clk_period;
Addr <= "1011111000001";
Trees_din <= "00000011000000000001111100000100";
wait for Clk_period;
Addr <= "1011111000010";
Trees_din <= "00000000001101110110000000110101";
wait for Clk_period;
Addr <= "1011111000011";
Trees_din <= "00000000001101110110000000110101";
wait for Clk_period;
Addr <= "1011111000100";
Trees_din <= "00000010000000000001100000000100";
wait for Clk_period;
Addr <= "1011111000101";
Trees_din <= "00000000000011010110000000110101";
wait for Clk_period;
Addr <= "1011111000110";
Trees_din <= "00000000000101000110000000110101";
wait for Clk_period;
Addr <= "1011111000111";
Trees_din <= "00000101000000000001011000001000";
wait for Clk_period;
Addr <= "1011111001000";
Trees_din <= "00000001000000000001101100000100";
wait for Clk_period;
Addr <= "1011111001001";
Trees_din <= "00000000000111000110000000110101";
wait for Clk_period;
Addr <= "1011111001010";
Trees_din <= "00000000001001000110000000110101";
wait for Clk_period;
Addr <= "1011111001011";
Trees_din <= "00000000000000000000111000000100";
wait for Clk_period;
Addr <= "1011111001100";
Trees_din <= "00000000001111110110000000110101";
wait for Clk_period;
Addr <= "1011111001101";
Trees_din <= "00000000010111000110000000110101";
wait for Clk_period;
Addr <= "1011111001110";
Trees_din <= "00000101000000000100111001000000";
wait for Clk_period;
Addr <= "1011111001111";
Trees_din <= "00000011000000000001000000100000";
wait for Clk_period;
Addr <= "1011111010000";
Trees_din <= "00000101000000000100000100010000";
wait for Clk_period;
Addr <= "1011111010001";
Trees_din <= "00000101000000000100010100001000";
wait for Clk_period;
Addr <= "1011111010010";
Trees_din <= "00000000000000000110001100000100";
wait for Clk_period;
Addr <= "1011111010011";
Trees_din <= "00000000000001000110000000110101";
wait for Clk_period;
Addr <= "1011111010100";
Trees_din <= "00000000010111100110000000110101";
wait for Clk_period;
Addr <= "1011111010101";
Trees_din <= "00000001000000000000111100000100";
wait for Clk_period;
Addr <= "1011111010110";
Trees_din <= "00000000010110110110000000110101";
wait for Clk_period;
Addr <= "1011111010111";
Trees_din <= "00000000001111010110000000110101";
wait for Clk_period;
Addr <= "1011111011000";
Trees_din <= "00000101000000000010101100001000";
wait for Clk_period;
Addr <= "1011111011001";
Trees_din <= "00000101000000000011010100000100";
wait for Clk_period;
Addr <= "1011111011010";
Trees_din <= "00000000000001100110000000110101";
wait for Clk_period;
Addr <= "1011111011011";
Trees_din <= "00000000000011000110000000110101";
wait for Clk_period;
Addr <= "1011111011100";
Trees_din <= "00000100000000000010100100000100";
wait for Clk_period;
Addr <= "1011111011101";
Trees_din <= "00000000010000000110000000110101";
wait for Clk_period;
Addr <= "1011111011110";
Trees_din <= "00000000000001000110000000110101";
wait for Clk_period;
Addr <= "1011111011111";
Trees_din <= "00000000000000000010011100010000";
wait for Clk_period;
Addr <= "1011111100000";
Trees_din <= "00000101000000000100010100001000";
wait for Clk_period;
Addr <= "1011111100001";
Trees_din <= "00000001000000000100000000000100";
wait for Clk_period;
Addr <= "1011111100010";
Trees_din <= "00000000001101100110000000110101";
wait for Clk_period;
Addr <= "1011111100011";
Trees_din <= "00000000000010010110000000110101";
wait for Clk_period;
Addr <= "1011111100100";
Trees_din <= "00000010000000000001000100000100";
wait for Clk_period;
Addr <= "1011111100101";
Trees_din <= "00000000000111110110000000110101";
wait for Clk_period;
Addr <= "1011111100110";
Trees_din <= "00000000010110010110000000110101";
wait for Clk_period;
Addr <= "1011111100111";
Trees_din <= "00000011000000000011110000001000";
wait for Clk_period;
Addr <= "1011111101000";
Trees_din <= "00000110000000000011111100000100";
wait for Clk_period;
Addr <= "1011111101001";
Trees_din <= "00000000010000100110000000110101";
wait for Clk_period;
Addr <= "1011111101010";
Trees_din <= "00000000010000100110000000110101";
wait for Clk_period;
Addr <= "1011111101011";
Trees_din <= "00000001000000000101110000000100";
wait for Clk_period;
Addr <= "1011111101100";
Trees_din <= "00000000001100000110000000110101";
wait for Clk_period;
Addr <= "1011111101101";
Trees_din <= "00000000010111000110000000110101";
wait for Clk_period;
Addr <= "1011111101110";
Trees_din <= "00000000000000000001100100100000";
wait for Clk_period;
Addr <= "1011111101111";
Trees_din <= "00000101000000000011110000010000";
wait for Clk_period;
Addr <= "1011111110000";
Trees_din <= "00000011000000000011001100001000";
wait for Clk_period;
Addr <= "1011111110001";
Trees_din <= "00000111000000000101100000000100";
wait for Clk_period;
Addr <= "1011111110010";
Trees_din <= "00000000001011010110000000110101";
wait for Clk_period;
Addr <= "1011111110011";
Trees_din <= "00000000010101100110000000110101";
wait for Clk_period;
Addr <= "1011111110100";
Trees_din <= "00000010000000000110001000000100";
wait for Clk_period;
Addr <= "1011111110101";
Trees_din <= "00000000000100100110000000110101";
wait for Clk_period;
Addr <= "1011111110110";
Trees_din <= "00000000001101010110000000110101";
wait for Clk_period;
Addr <= "1011111110111";
Trees_din <= "00000101000000000010000100001000";
wait for Clk_period;
Addr <= "1011111111000";
Trees_din <= "00000100000000000011000000000100";
wait for Clk_period;
Addr <= "1011111111001";
Trees_din <= "00000000000111010110000000110101";
wait for Clk_period;
Addr <= "1011111111010";
Trees_din <= "00000000010101110110000000110101";
wait for Clk_period;
Addr <= "1011111111011";
Trees_din <= "00000001000000000110000000000100";
wait for Clk_period;
Addr <= "1011111111100";
Trees_din <= "00000000010010000110000000110101";
wait for Clk_period;
Addr <= "1011111111101";
Trees_din <= "00000000010100100110000000110101";
wait for Clk_period;
Addr <= "1011111111110";
Trees_din <= "00000010000000000001001100010000";
wait for Clk_period;
Addr <= "1011111111111";
Trees_din <= "00000110000000000000100000001000";
wait for Clk_period;
Addr <= "1100000000000";
Trees_din <= "00000010000000000110001100000100";
wait for Clk_period;
Addr <= "1100000000001";
Trees_din <= "00000000000111100110000000110101";
wait for Clk_period;
Addr <= "1100000000010";
Trees_din <= "00000000000010100110000000110101";
wait for Clk_period;
Addr <= "1100000000011";
Trees_din <= "00000111000000000101000100000100";
wait for Clk_period;
Addr <= "1100000000100";
Trees_din <= "00000000001000110110000000110101";
wait for Clk_period;
Addr <= "1100000000101";
Trees_din <= "00000000001100010110000000110101";
wait for Clk_period;
Addr <= "1100000000110";
Trees_din <= "00000111000000000011110000001000";
wait for Clk_period;
Addr <= "1100000000111";
Trees_din <= "00000111000000000101100100000100";
wait for Clk_period;
Addr <= "1100000001000";
Trees_din <= "00000000010101110110000000110101";
wait for Clk_period;
Addr <= "1100000001001";
Trees_din <= "00000000000011010110000000110101";
wait for Clk_period;
Addr <= "1100000001010";
Trees_din <= "00000101000000000011111100000100";
wait for Clk_period;
Addr <= "1100000001011";
Trees_din <= "00000000001111100110000000110101";
wait for Clk_period;
Addr <= "1100000001100";
Trees_din <= "00000000000111000110000000110101";
wait for Clk_period;



----------tree 48-------------------

Addr <= "1100000001101";
Trees_din <= "00000011000000000100010110000000";
wait for Clk_period;
Addr <= "1100000001110";
Trees_din <= "00000001000000000100100101000000";
wait for Clk_period;
Addr <= "1100000001111";
Trees_din <= "00000011000000000011100100100000";
wait for Clk_period;
Addr <= "1100000010000";
Trees_din <= "00000001000000000010100100010000";
wait for Clk_period;
Addr <= "1100000010001";
Trees_din <= "00000101000000000101011100001000";
wait for Clk_period;
Addr <= "1100000010010";
Trees_din <= "00000100000000000011110000000100";
wait for Clk_period;
Addr <= "1100000010011";
Trees_din <= "00000000000010100110001000110001";
wait for Clk_period;
Addr <= "1100000010100";
Trees_din <= "00000000000101000110001000110001";
wait for Clk_period;
Addr <= "1100000010101";
Trees_din <= "00000100000000000010010000000100";
wait for Clk_period;
Addr <= "1100000010110";
Trees_din <= "00000000000000100110001000110001";
wait for Clk_period;
Addr <= "1100000010111";
Trees_din <= "00000000001110000110001000110001";
wait for Clk_period;
Addr <= "1100000011000";
Trees_din <= "00000011000000000010000000001000";
wait for Clk_period;
Addr <= "1100000011001";
Trees_din <= "00000010000000000000000000000100";
wait for Clk_period;
Addr <= "1100000011010";
Trees_din <= "00000000001100110110001000110001";
wait for Clk_period;
Addr <= "1100000011011";
Trees_din <= "00000000001101010110001000110001";
wait for Clk_period;
Addr <= "1100000011100";
Trees_din <= "00000110000000000001101000000100";
wait for Clk_period;
Addr <= "1100000011101";
Trees_din <= "00000000010110100110001000110001";
wait for Clk_period;
Addr <= "1100000011110";
Trees_din <= "00000000000001010110001000110001";
wait for Clk_period;
Addr <= "1100000011111";
Trees_din <= "00000011000000000011001000010000";
wait for Clk_period;
Addr <= "1100000100000";
Trees_din <= "00000001000000000011001000001000";
wait for Clk_period;
Addr <= "1100000100001";
Trees_din <= "00000000000000000001000000000100";
wait for Clk_period;
Addr <= "1100000100010";
Trees_din <= "00000000000011010110001000110001";
wait for Clk_period;
Addr <= "1100000100011";
Trees_din <= "00000000000000100110001000110001";
wait for Clk_period;
Addr <= "1100000100100";
Trees_din <= "00000100000000000011011100000100";
wait for Clk_period;
Addr <= "1100000100101";
Trees_din <= "00000000010111110110001000110001";
wait for Clk_period;
Addr <= "1100000100110";
Trees_din <= "00000000000001000110001000110001";
wait for Clk_period;
Addr <= "1100000100111";
Trees_din <= "00000111000000000001011100001000";
wait for Clk_period;
Addr <= "1100000101000";
Trees_din <= "00000111000000000001000100000100";
wait for Clk_period;
Addr <= "1100000101001";
Trees_din <= "00000000000100010110001000110001";
wait for Clk_period;
Addr <= "1100000101010";
Trees_din <= "00000000000111100110001000110001";
wait for Clk_period;
Addr <= "1100000101011";
Trees_din <= "00000101000000000000010000000100";
wait for Clk_period;
Addr <= "1100000101100";
Trees_din <= "00000000001110000110001000110001";
wait for Clk_period;
Addr <= "1100000101101";
Trees_din <= "00000000000010000110001000110001";
wait for Clk_period;
Addr <= "1100000101110";
Trees_din <= "00000100000000000001001100100000";
wait for Clk_period;
Addr <= "1100000101111";
Trees_din <= "00000101000000000100111000010000";
wait for Clk_period;
Addr <= "1100000110000";
Trees_din <= "00000001000000000100010100001000";
wait for Clk_period;
Addr <= "1100000110001";
Trees_din <= "00000001000000000100011100000100";
wait for Clk_period;
Addr <= "1100000110010";
Trees_din <= "00000000000001110110001000110001";
wait for Clk_period;
Addr <= "1100000110011";
Trees_din <= "00000000010011010110001000110001";
wait for Clk_period;
Addr <= "1100000110100";
Trees_din <= "00000001000000000010101000000100";
wait for Clk_period;
Addr <= "1100000110101";
Trees_din <= "00000000000000110110001000110001";
wait for Clk_period;
Addr <= "1100000110110";
Trees_din <= "00000000000011000110001000110001";
wait for Clk_period;
Addr <= "1100000110111";
Trees_din <= "00000001000000000010011000001000";
wait for Clk_period;
Addr <= "1100000111000";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "1100000111001";
Trees_din <= "00000000010101000110001000110001";
wait for Clk_period;
Addr <= "1100000111010";
Trees_din <= "00000000000010000110001000110001";
wait for Clk_period;
Addr <= "1100000111011";
Trees_din <= "00000010000000000010111100000100";
wait for Clk_period;
Addr <= "1100000111100";
Trees_din <= "00000000001101110110001000110001";
wait for Clk_period;
Addr <= "1100000111101";
Trees_din <= "00000000000111110110001000110001";
wait for Clk_period;
Addr <= "1100000111110";
Trees_din <= "00000110000000000011101100010000";
wait for Clk_period;
Addr <= "1100000111111";
Trees_din <= "00000001000000000010101100001000";
wait for Clk_period;
Addr <= "1100001000000";
Trees_din <= "00000001000000000101110000000100";
wait for Clk_period;
Addr <= "1100001000001";
Trees_din <= "00000000001100010110001000110001";
wait for Clk_period;
Addr <= "1100001000010";
Trees_din <= "00000000010001010110001000110001";
wait for Clk_period;
Addr <= "1100001000011";
Trees_din <= "00000000000000000001100000000100";
wait for Clk_period;
Addr <= "1100001000100";
Trees_din <= "00000000000000100110001000110001";
wait for Clk_period;
Addr <= "1100001000101";
Trees_din <= "00000000010001100110001000110001";
wait for Clk_period;
Addr <= "1100001000110";
Trees_din <= "00000100000000000010100100001000";
wait for Clk_period;
Addr <= "1100001000111";
Trees_din <= "00000010000000000101000100000100";
wait for Clk_period;
Addr <= "1100001001000";
Trees_din <= "00000000010100010110001000110001";
wait for Clk_period;
Addr <= "1100001001001";
Trees_din <= "00000000001110000110001000110001";
wait for Clk_period;
Addr <= "1100001001010";
Trees_din <= "00000000000000000100001100000100";
wait for Clk_period;
Addr <= "1100001001011";
Trees_din <= "00000000001000000110001000110001";
wait for Clk_period;
Addr <= "1100001001100";
Trees_din <= "00000000010001000110001000110001";
wait for Clk_period;
Addr <= "1100001001101";
Trees_din <= "00000001000000000010111001000000";
wait for Clk_period;
Addr <= "1100001001110";
Trees_din <= "00000011000000000010100100100000";
wait for Clk_period;
Addr <= "1100001001111";
Trees_din <= "00000011000000000101110100010000";
wait for Clk_period;
Addr <= "1100001010000";
Trees_din <= "00000100000000000110010000001000";
wait for Clk_period;
Addr <= "1100001010001";
Trees_din <= "00000000000000000100000000000100";
wait for Clk_period;
Addr <= "1100001010010";
Trees_din <= "00000000010010000110001000110001";
wait for Clk_period;
Addr <= "1100001010011";
Trees_din <= "00000000010101100110001000110001";
wait for Clk_period;
Addr <= "1100001010100";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "1100001010101";
Trees_din <= "00000000001010000110001000110001";
wait for Clk_period;
Addr <= "1100001010110";
Trees_din <= "00000000000000110110001000110001";
wait for Clk_period;
Addr <= "1100001010111";
Trees_din <= "00000011000000000010010000001000";
wait for Clk_period;
Addr <= "1100001011000";
Trees_din <= "00000110000000000011010000000100";
wait for Clk_period;
Addr <= "1100001011001";
Trees_din <= "00000000010111100110001000110001";
wait for Clk_period;
Addr <= "1100001011010";
Trees_din <= "00000000001000000110001000110001";
wait for Clk_period;
Addr <= "1100001011011";
Trees_din <= "00000000000000000001010000000100";
wait for Clk_period;
Addr <= "1100001011100";
Trees_din <= "00000000001001010110001000110001";
wait for Clk_period;
Addr <= "1100001011101";
Trees_din <= "00000000001010100110001000110001";
wait for Clk_period;
Addr <= "1100001011110";
Trees_din <= "00000101000000000011011000010000";
wait for Clk_period;
Addr <= "1100001011111";
Trees_din <= "00000010000000000100001100001000";
wait for Clk_period;
Addr <= "1100001100000";
Trees_din <= "00000111000000000000001100000100";
wait for Clk_period;
Addr <= "1100001100001";
Trees_din <= "00000000001110010110001000110001";
wait for Clk_period;
Addr <= "1100001100010";
Trees_din <= "00000000011000000110001000110001";
wait for Clk_period;
Addr <= "1100001100011";
Trees_din <= "00000111000000000001000000000100";
wait for Clk_period;
Addr <= "1100001100100";
Trees_din <= "00000000001100110110001000110001";
wait for Clk_period;
Addr <= "1100001100101";
Trees_din <= "00000000010111110110001000110001";
wait for Clk_period;
Addr <= "1100001100110";
Trees_din <= "00000111000000000110010000001000";
wait for Clk_period;
Addr <= "1100001100111";
Trees_din <= "00000000000000000100010100000100";
wait for Clk_period;
Addr <= "1100001101000";
Trees_din <= "00000000010100000110001000110001";
wait for Clk_period;
Addr <= "1100001101001";
Trees_din <= "00000000010000110110001000110001";
wait for Clk_period;
Addr <= "1100001101010";
Trees_din <= "00000000000000000011101000000100";
wait for Clk_period;
Addr <= "1100001101011";
Trees_din <= "00000000000000110110001000110001";
wait for Clk_period;
Addr <= "1100001101100";
Trees_din <= "00000000000110110110001000110001";
wait for Clk_period;
Addr <= "1100001101101";
Trees_din <= "00000111000000000011110100100000";
wait for Clk_period;
Addr <= "1100001101110";
Trees_din <= "00000010000000000000110000010000";
wait for Clk_period;
Addr <= "1100001101111";
Trees_din <= "00000000000000000011000000001000";
wait for Clk_period;
Addr <= "1100001110000";
Trees_din <= "00000111000000000101000100000100";
wait for Clk_period;
Addr <= "1100001110001";
Trees_din <= "00000000000000100110001000110001";
wait for Clk_period;
Addr <= "1100001110010";
Trees_din <= "00000000010110000110001000110001";
wait for Clk_period;
Addr <= "1100001110011";
Trees_din <= "00000001000000000101110100000100";
wait for Clk_period;
Addr <= "1100001110100";
Trees_din <= "00000000001011010110001000110001";
wait for Clk_period;
Addr <= "1100001110101";
Trees_din <= "00000000000111010110001000110001";
wait for Clk_period;
Addr <= "1100001110110";
Trees_din <= "00000010000000000011111000001000";
wait for Clk_period;
Addr <= "1100001110111";
Trees_din <= "00000000000000000001000000000100";
wait for Clk_period;
Addr <= "1100001111000";
Trees_din <= "00000000010110000110001000110001";
wait for Clk_period;
Addr <= "1100001111001";
Trees_din <= "00000000001101100110001000110001";
wait for Clk_period;
Addr <= "1100001111010";
Trees_din <= "00000010000000000100010100000100";
wait for Clk_period;
Addr <= "1100001111011";
Trees_din <= "00000000010101000110001000110001";
wait for Clk_period;
Addr <= "1100001111100";
Trees_din <= "00000000000100100110001000110001";
wait for Clk_period;
Addr <= "1100001111101";
Trees_din <= "00000101000000000000110100010000";
wait for Clk_period;
Addr <= "1100001111110";
Trees_din <= "00000011000000000001001100001000";
wait for Clk_period;
Addr <= "1100001111111";
Trees_din <= "00000100000000000010000100000100";
wait for Clk_period;
Addr <= "1100010000000";
Trees_din <= "00000000010000100110001000110001";
wait for Clk_period;
Addr <= "1100010000001";
Trees_din <= "00000000000011110110001000110001";
wait for Clk_period;
Addr <= "1100010000010";
Trees_din <= "00000110000000000101101100000100";
wait for Clk_period;
Addr <= "1100010000011";
Trees_din <= "00000000000000000110001000110001";
wait for Clk_period;
Addr <= "1100010000100";
Trees_din <= "00000000001101000110001000110001";
wait for Clk_period;
Addr <= "1100010000101";
Trees_din <= "00000101000000000100010000001000";
wait for Clk_period;
Addr <= "1100010000110";
Trees_din <= "00000110000000000000001100000100";
wait for Clk_period;
Addr <= "1100010000111";
Trees_din <= "00000000001111000110001000110001";
wait for Clk_period;
Addr <= "1100010001000";
Trees_din <= "00000000001001000110001000110001";
wait for Clk_period;
Addr <= "1100010001001";
Trees_din <= "00000011000000000000111100000100";
wait for Clk_period;
Addr <= "1100010001010";
Trees_din <= "00000000000001010110001000110001";
wait for Clk_period;
Addr <= "1100010001011";
Trees_din <= "00000000010111110110001000110001";
wait for Clk_period;



----------tree 49-------------------

Addr <= "1100010001100";
Trees_din <= "00000000000000000101011010000000";
wait for Clk_period;
Addr <= "1100010001101";
Trees_din <= "00000101000000000000011001000000";
wait for Clk_period;
Addr <= "1100010001110";
Trees_din <= "00000100000000000001111100100000";
wait for Clk_period;
Addr <= "1100010001111";
Trees_din <= "00000110000000000001110000010000";
wait for Clk_period;
Addr <= "1100010010000";
Trees_din <= "00000101000000000011011100001000";
wait for Clk_period;
Addr <= "1100010010001";
Trees_din <= "00000011000000000001100000000100";
wait for Clk_period;
Addr <= "1100010010010";
Trees_din <= "00000000001000100110010000101111";
wait for Clk_period;
Addr <= "1100010010011";
Trees_din <= "00000000010011010110010000101111";
wait for Clk_period;
Addr <= "1100010010100";
Trees_din <= "00000111000000000100100000000100";
wait for Clk_period;
Addr <= "1100010010101";
Trees_din <= "00000000000001010110010000101111";
wait for Clk_period;
Addr <= "1100010010110";
Trees_din <= "00000000010001000110010000101111";
wait for Clk_period;
Addr <= "1100010010111";
Trees_din <= "00000100000000000000011100001000";
wait for Clk_period;
Addr <= "1100010011000";
Trees_din <= "00000111000000000100111100000100";
wait for Clk_period;
Addr <= "1100010011001";
Trees_din <= "00000000000010000110010000101111";
wait for Clk_period;
Addr <= "1100010011010";
Trees_din <= "00000000000001010110010000101111";
wait for Clk_period;
Addr <= "1100010011011";
Trees_din <= "00000111000000000000010100000100";
wait for Clk_period;
Addr <= "1100010011100";
Trees_din <= "00000000010000100110010000101111";
wait for Clk_period;
Addr <= "1100010011101";
Trees_din <= "00000000010010100110010000101111";
wait for Clk_period;
Addr <= "1100010011110";
Trees_din <= "00000010000000000101100000010000";
wait for Clk_period;
Addr <= "1100010011111";
Trees_din <= "00000110000000000011001100001000";
wait for Clk_period;
Addr <= "1100010100000";
Trees_din <= "00000110000000000101000100000100";
wait for Clk_period;
Addr <= "1100010100001";
Trees_din <= "00000000000100000110010000101111";
wait for Clk_period;
Addr <= "1100010100010";
Trees_din <= "00000000001001110110010000101111";
wait for Clk_period;
Addr <= "1100010100011";
Trees_din <= "00000011000000000101001100000100";
wait for Clk_period;
Addr <= "1100010100100";
Trees_din <= "00000000010111110110010000101111";
wait for Clk_period;
Addr <= "1100010100101";
Trees_din <= "00000000001000010110010000101111";
wait for Clk_period;
Addr <= "1100010100110";
Trees_din <= "00000101000000000110010000001000";
wait for Clk_period;
Addr <= "1100010100111";
Trees_din <= "00000011000000000010110000000100";
wait for Clk_period;
Addr <= "1100010101000";
Trees_din <= "00000000010101010110010000101111";
wait for Clk_period;
Addr <= "1100010101001";
Trees_din <= "00000000010010110110010000101111";
wait for Clk_period;
Addr <= "1100010101010";
Trees_din <= "00000100000000000100111000000100";
wait for Clk_period;
Addr <= "1100010101011";
Trees_din <= "00000000000101110110010000101111";
wait for Clk_period;
Addr <= "1100010101100";
Trees_din <= "00000000001000000110010000101111";
wait for Clk_period;
Addr <= "1100010101101";
Trees_din <= "00000101000000000110010000100000";
wait for Clk_period;
Addr <= "1100010101110";
Trees_din <= "00000101000000000010001100010000";
wait for Clk_period;
Addr <= "1100010101111";
Trees_din <= "00000000000000000100010000001000";
wait for Clk_period;
Addr <= "1100010110000";
Trees_din <= "00000111000000000001001000000100";
wait for Clk_period;
Addr <= "1100010110001";
Trees_din <= "00000000000111000110010000101111";
wait for Clk_period;
Addr <= "1100010110010";
Trees_din <= "00000000000101010110010000101111";
wait for Clk_period;
Addr <= "1100010110011";
Trees_din <= "00000011000000000000100100000100";
wait for Clk_period;
Addr <= "1100010110100";
Trees_din <= "00000000001101000110010000101111";
wait for Clk_period;
Addr <= "1100010110101";
Trees_din <= "00000000010001000110010000101111";
wait for Clk_period;
Addr <= "1100010110110";
Trees_din <= "00000100000000000110001100001000";
wait for Clk_period;
Addr <= "1100010110111";
Trees_din <= "00000110000000000000110100000100";
wait for Clk_period;
Addr <= "1100010111000";
Trees_din <= "00000000010010110110010000101111";
wait for Clk_period;
Addr <= "1100010111001";
Trees_din <= "00000000010111100110010000101111";
wait for Clk_period;
Addr <= "1100010111010";
Trees_din <= "00000010000000000000010100000100";
wait for Clk_period;
Addr <= "1100010111011";
Trees_din <= "00000000000100000110010000101111";
wait for Clk_period;
Addr <= "1100010111100";
Trees_din <= "00000000001010110110010000101111";
wait for Clk_period;
Addr <= "1100010111101";
Trees_din <= "00000000000000000101110100010000";
wait for Clk_period;
Addr <= "1100010111110";
Trees_din <= "00000001000000000010000100001000";
wait for Clk_period;
Addr <= "1100010111111";
Trees_din <= "00000110000000000101011100000100";
wait for Clk_period;
Addr <= "1100011000000";
Trees_din <= "00000000001110010110010000101111";
wait for Clk_period;
Addr <= "1100011000001";
Trees_din <= "00000000000100100110010000101111";
wait for Clk_period;
Addr <= "1100011000010";
Trees_din <= "00000111000000000000101000000100";
wait for Clk_period;
Addr <= "1100011000011";
Trees_din <= "00000000001101010110010000101111";
wait for Clk_period;
Addr <= "1100011000100";
Trees_din <= "00000000000000100110010000101111";
wait for Clk_period;
Addr <= "1100011000101";
Trees_din <= "00000011000000000101011100001000";
wait for Clk_period;
Addr <= "1100011000110";
Trees_din <= "00000010000000000011100000000100";
wait for Clk_period;
Addr <= "1100011000111";
Trees_din <= "00000000001001000110010000101111";
wait for Clk_period;
Addr <= "1100011001000";
Trees_din <= "00000000000100110110010000101111";
wait for Clk_period;
Addr <= "1100011001001";
Trees_din <= "00000001000000000001010100000100";
wait for Clk_period;
Addr <= "1100011001010";
Trees_din <= "00000000010100110110010000101111";
wait for Clk_period;
Addr <= "1100011001011";
Trees_din <= "00000000010001100110010000101111";
wait for Clk_period;
Addr <= "1100011001100";
Trees_din <= "00000110000000000001001001000000";
wait for Clk_period;
Addr <= "1100011001101";
Trees_din <= "00000111000000000001101000100000";
wait for Clk_period;
Addr <= "1100011001110";
Trees_din <= "00000111000000000010101100010000";
wait for Clk_period;
Addr <= "1100011001111";
Trees_din <= "00000010000000000010011100001000";
wait for Clk_period;
Addr <= "1100011010000";
Trees_din <= "00000001000000000011000000000100";
wait for Clk_period;
Addr <= "1100011010001";
Trees_din <= "00000000000001100110010000101111";
wait for Clk_period;
Addr <= "1100011010010";
Trees_din <= "00000000010110100110010000101111";
wait for Clk_period;
Addr <= "1100011010011";
Trees_din <= "00000111000000000110000100000100";
wait for Clk_period;
Addr <= "1100011010100";
Trees_din <= "00000000010101110110010000101111";
wait for Clk_period;
Addr <= "1100011010101";
Trees_din <= "00000000000001010110010000101111";
wait for Clk_period;
Addr <= "1100011010110";
Trees_din <= "00000111000000000010101000001000";
wait for Clk_period;
Addr <= "1100011010111";
Trees_din <= "00000100000000000110000000000100";
wait for Clk_period;
Addr <= "1100011011000";
Trees_din <= "00000000010011110110010000101111";
wait for Clk_period;
Addr <= "1100011011001";
Trees_din <= "00000000000000100110010000101111";
wait for Clk_period;
Addr <= "1100011011010";
Trees_din <= "00000100000000000001010000000100";
wait for Clk_period;
Addr <= "1100011011011";
Trees_din <= "00000000000011000110010000101111";
wait for Clk_period;
Addr <= "1100011011100";
Trees_din <= "00000000010001010110010000101111";
wait for Clk_period;
Addr <= "1100011011101";
Trees_din <= "00000101000000000100100100010000";
wait for Clk_period;
Addr <= "1100011011110";
Trees_din <= "00000110000000000001111000001000";
wait for Clk_period;
Addr <= "1100011011111";
Trees_din <= "00000100000000000101001000000100";
wait for Clk_period;
Addr <= "1100011100000";
Trees_din <= "00000000010011010110010000101111";
wait for Clk_period;
Addr <= "1100011100001";
Trees_din <= "00000000000100100110010000101111";
wait for Clk_period;
Addr <= "1100011100010";
Trees_din <= "00000100000000000001110100000100";
wait for Clk_period;
Addr <= "1100011100011";
Trees_din <= "00000000000100010110010000101111";
wait for Clk_period;
Addr <= "1100011100100";
Trees_din <= "00000000001111100110010000101111";
wait for Clk_period;
Addr <= "1100011100101";
Trees_din <= "00000010000000000100000000001000";
wait for Clk_period;
Addr <= "1100011100110";
Trees_din <= "00000101000000000010010100000100";
wait for Clk_period;
Addr <= "1100011100111";
Trees_din <= "00000000001110110110010000101111";
wait for Clk_period;
Addr <= "1100011101000";
Trees_din <= "00000000010101110110010000101111";
wait for Clk_period;
Addr <= "1100011101001";
Trees_din <= "00000001000000000001110100000100";
wait for Clk_period;
Addr <= "1100011101010";
Trees_din <= "00000000010000100110010000101111";
wait for Clk_period;
Addr <= "1100011101011";
Trees_din <= "00000000010000000110010000101111";
wait for Clk_period;
Addr <= "1100011101100";
Trees_din <= "00000010000000000100100000100000";
wait for Clk_period;
Addr <= "1100011101101";
Trees_din <= "00000011000000000011000100010000";
wait for Clk_period;
Addr <= "1100011101110";
Trees_din <= "00000001000000000011111100001000";
wait for Clk_period;
Addr <= "1100011101111";
Trees_din <= "00000111000000000011110100000100";
wait for Clk_period;
Addr <= "1100011110000";
Trees_din <= "00000000001110010110010000101111";
wait for Clk_period;
Addr <= "1100011110001";
Trees_din <= "00000000010100000110010000101111";
wait for Clk_period;
Addr <= "1100011110010";
Trees_din <= "00000010000000000000011000000100";
wait for Clk_period;
Addr <= "1100011110011";
Trees_din <= "00000000001110010110010000101111";
wait for Clk_period;
Addr <= "1100011110100";
Trees_din <= "00000000000100110110010000101111";
wait for Clk_period;
Addr <= "1100011110101";
Trees_din <= "00000001000000000001001100001000";
wait for Clk_period;
Addr <= "1100011110110";
Trees_din <= "00000011000000000011111000000100";
wait for Clk_period;
Addr <= "1100011110111";
Trees_din <= "00000000010011100110010000101111";
wait for Clk_period;
Addr <= "1100011111000";
Trees_din <= "00000000010101010110010000101111";
wait for Clk_period;
Addr <= "1100011111001";
Trees_din <= "00000110000000000101101100000100";
wait for Clk_period;
Addr <= "1100011111010";
Trees_din <= "00000000010011010110010000101111";
wait for Clk_period;
Addr <= "1100011111011";
Trees_din <= "00000000010110000110010000101111";
wait for Clk_period;
Addr <= "1100011111100";
Trees_din <= "00000101000000000000100000010000";
wait for Clk_period;
Addr <= "1100011111101";
Trees_din <= "00000011000000000010011000001000";
wait for Clk_period;
Addr <= "1100011111110";
Trees_din <= "00000010000000000000100000000100";
wait for Clk_period;
Addr <= "1100011111111";
Trees_din <= "00000000001101000110010000101111";
wait for Clk_period;
Addr <= "1100100000000";
Trees_din <= "00000000000001110110010000101111";
wait for Clk_period;
Addr <= "1100100000001";
Trees_din <= "00000101000000000011001100000100";
wait for Clk_period;
Addr <= "1100100000010";
Trees_din <= "00000000000111010110010000101111";
wait for Clk_period;
Addr <= "1100100000011";
Trees_din <= "00000000010101110110010000101111";
wait for Clk_period;
Addr <= "1100100000100";
Trees_din <= "00000100000000000001111100001000";
wait for Clk_period;
Addr <= "1100100000101";
Trees_din <= "00000100000000000101000000000100";
wait for Clk_period;
Addr <= "1100100000110";
Trees_din <= "00000000010001010110010000101111";
wait for Clk_period;
Addr <= "1100100000111";
Trees_din <= "00000000000011000110010000101111";
wait for Clk_period;
Addr <= "1100100001000";
Trees_din <= "00000110000000000001010100000100";
wait for Clk_period;
Addr <= "1100100001001";
Trees_din <= "00000000001011100110010000101111";
wait for Clk_period;
Addr <= "1100100001010";
Trees_din <= "00000000010000010110010000101111";
wait for Clk_period;



----------tree 50-------------------

Addr <= "1100100001011";
Trees_din <= "00000101000000000101000110000000";
wait for Clk_period;
Addr <= "1100100001100";
Trees_din <= "00000111000000000010010001000000";
wait for Clk_period;
Addr <= "1100100001101";
Trees_din <= "00000110000000000101110100100000";
wait for Clk_period;
Addr <= "1100100001110";
Trees_din <= "00000001000000000001111100010000";
wait for Clk_period;
Addr <= "1100100001111";
Trees_din <= "00000101000000000011000100001000";
wait for Clk_period;
Addr <= "1100100010000";
Trees_din <= "00000110000000000101101100000100";
wait for Clk_period;
Addr <= "1100100010001";
Trees_din <= "00000000000111010110011000101001";
wait for Clk_period;
Addr <= "1100100010010";
Trees_din <= "00000000001001010110011000101001";
wait for Clk_period;
Addr <= "1100100010011";
Trees_din <= "00000101000000000100001100000100";
wait for Clk_period;
Addr <= "1100100010100";
Trees_din <= "00000000010111100110011000101001";
wait for Clk_period;
Addr <= "1100100010101";
Trees_din <= "00000000010110100110011000101001";
wait for Clk_period;
Addr <= "1100100010110";
Trees_din <= "00000010000000000100101000001000";
wait for Clk_period;
Addr <= "1100100010111";
Trees_din <= "00000111000000000010010100000100";
wait for Clk_period;
Addr <= "1100100011000";
Trees_din <= "00000000010000110110011000101001";
wait for Clk_period;
Addr <= "1100100011001";
Trees_din <= "00000000000010110110011000101001";
wait for Clk_period;
Addr <= "1100100011010";
Trees_din <= "00000010000000000000001100000100";
wait for Clk_period;
Addr <= "1100100011011";
Trees_din <= "00000000001001110110011000101001";
wait for Clk_period;
Addr <= "1100100011100";
Trees_din <= "00000000001011110110011000101001";
wait for Clk_period;
Addr <= "1100100011101";
Trees_din <= "00000001000000000011110000010000";
wait for Clk_period;
Addr <= "1100100011110";
Trees_din <= "00000001000000000101101100001000";
wait for Clk_period;
Addr <= "1100100011111";
Trees_din <= "00000111000000000101110000000100";
wait for Clk_period;
Addr <= "1100100100000";
Trees_din <= "00000000010100010110011000101001";
wait for Clk_period;
Addr <= "1100100100001";
Trees_din <= "00000000010111100110011000101001";
wait for Clk_period;
Addr <= "1100100100010";
Trees_din <= "00000011000000000101000100000100";
wait for Clk_period;
Addr <= "1100100100011";
Trees_din <= "00000000000000000110011000101001";
wait for Clk_period;
Addr <= "1100100100100";
Trees_din <= "00000000000001100110011000101001";
wait for Clk_period;
Addr <= "1100100100101";
Trees_din <= "00000010000000000011000100001000";
wait for Clk_period;
Addr <= "1100100100110";
Trees_din <= "00000101000000000100010000000100";
wait for Clk_period;
Addr <= "1100100100111";
Trees_din <= "00000000001100100110011000101001";
wait for Clk_period;
Addr <= "1100100101000";
Trees_din <= "00000000001100100110011000101001";
wait for Clk_period;
Addr <= "1100100101001";
Trees_din <= "00000100000000000101101100000100";
wait for Clk_period;
Addr <= "1100100101010";
Trees_din <= "00000000001011100110011000101001";
wait for Clk_period;
Addr <= "1100100101011";
Trees_din <= "00000000010101010110011000101001";
wait for Clk_period;
Addr <= "1100100101100";
Trees_din <= "00000100000000000101110000100000";
wait for Clk_period;
Addr <= "1100100101101";
Trees_din <= "00000110000000000010011000010000";
wait for Clk_period;
Addr <= "1100100101110";
Trees_din <= "00000000000000000101100000001000";
wait for Clk_period;
Addr <= "1100100101111";
Trees_din <= "00000001000000000000010100000100";
wait for Clk_period;
Addr <= "1100100110000";
Trees_din <= "00000000010001100110011000101001";
wait for Clk_period;
Addr <= "1100100110001";
Trees_din <= "00000000000110110110011000101001";
wait for Clk_period;
Addr <= "1100100110010";
Trees_din <= "00000010000000000010101000000100";
wait for Clk_period;
Addr <= "1100100110011";
Trees_din <= "00000000010011010110011000101001";
wait for Clk_period;
Addr <= "1100100110100";
Trees_din <= "00000000010011100110011000101001";
wait for Clk_period;
Addr <= "1100100110101";
Trees_din <= "00000010000000000101010000001000";
wait for Clk_period;
Addr <= "1100100110110";
Trees_din <= "00000000000000000011011000000100";
wait for Clk_period;
Addr <= "1100100110111";
Trees_din <= "00000000001111110110011000101001";
wait for Clk_period;
Addr <= "1100100111000";
Trees_din <= "00000000001110000110011000101001";
wait for Clk_period;
Addr <= "1100100111001";
Trees_din <= "00000011000000000100110100000100";
wait for Clk_period;
Addr <= "1100100111010";
Trees_din <= "00000000010011010110011000101001";
wait for Clk_period;
Addr <= "1100100111011";
Trees_din <= "00000000001001110110011000101001";
wait for Clk_period;
Addr <= "1100100111100";
Trees_din <= "00000000000000000011000000010000";
wait for Clk_period;
Addr <= "1100100111101";
Trees_din <= "00000001000000000110000000001000";
wait for Clk_period;
Addr <= "1100100111110";
Trees_din <= "00000001000000000101010000000100";
wait for Clk_period;
Addr <= "1100100111111";
Trees_din <= "00000000001010010110011000101001";
wait for Clk_period;
Addr <= "1100101000000";
Trees_din <= "00000000010100000110011000101001";
wait for Clk_period;
Addr <= "1100101000001";
Trees_din <= "00000101000000000011001100000100";
wait for Clk_period;
Addr <= "1100101000010";
Trees_din <= "00000000011001000110011000101001";
wait for Clk_period;
Addr <= "1100101000011";
Trees_din <= "00000000010110000110011000101001";
wait for Clk_period;
Addr <= "1100101000100";
Trees_din <= "00000101000000000001100000001000";
wait for Clk_period;
Addr <= "1100101000101";
Trees_din <= "00000100000000000110000100000100";
wait for Clk_period;
Addr <= "1100101000110";
Trees_din <= "00000000011000110110011000101001";
wait for Clk_period;
Addr <= "1100101000111";
Trees_din <= "00000000000111010110011000101001";
wait for Clk_period;
Addr <= "1100101001000";
Trees_din <= "00000001000000000100011100000100";
wait for Clk_period;
Addr <= "1100101001001";
Trees_din <= "00000000001100000110011000101001";
wait for Clk_period;
Addr <= "1100101001010";
Trees_din <= "00000000000101100110011000101001";
wait for Clk_period;
Addr <= "1100101001011";
Trees_din <= "00000101000000000101110001000000";
wait for Clk_period;
Addr <= "1100101001100";
Trees_din <= "00000001000000000100110100100000";
wait for Clk_period;
Addr <= "1100101001101";
Trees_din <= "00000110000000000000000100010000";
wait for Clk_period;
Addr <= "1100101001110";
Trees_din <= "00000110000000000100001100001000";
wait for Clk_period;
Addr <= "1100101001111";
Trees_din <= "00000010000000000010110100000100";
wait for Clk_period;
Addr <= "1100101010000";
Trees_din <= "00000000000010100110011000101001";
wait for Clk_period;
Addr <= "1100101010001";
Trees_din <= "00000000011000000110011000101001";
wait for Clk_period;
Addr <= "1100101010010";
Trees_din <= "00000000000000000101010000000100";
wait for Clk_period;
Addr <= "1100101010011";
Trees_din <= "00000000010100110110011000101001";
wait for Clk_period;
Addr <= "1100101010100";
Trees_din <= "00000000000010110110011000101001";
wait for Clk_period;
Addr <= "1100101010101";
Trees_din <= "00000111000000000100000000001000";
wait for Clk_period;
Addr <= "1100101010110";
Trees_din <= "00000101000000000011100000000100";
wait for Clk_period;
Addr <= "1100101010111";
Trees_din <= "00000000010011110110011000101001";
wait for Clk_period;
Addr <= "1100101011000";
Trees_din <= "00000000010110110110011000101001";
wait for Clk_period;
Addr <= "1100101011001";
Trees_din <= "00000110000000000010110000000100";
wait for Clk_period;
Addr <= "1100101011010";
Trees_din <= "00000000001010010110011000101001";
wait for Clk_period;
Addr <= "1100101011011";
Trees_din <= "00000000010111110110011000101001";
wait for Clk_period;
Addr <= "1100101011100";
Trees_din <= "00000101000000000101110000010000";
wait for Clk_period;
Addr <= "1100101011101";
Trees_din <= "00000001000000000010011100001000";
wait for Clk_period;
Addr <= "1100101011110";
Trees_din <= "00000011000000000000011000000100";
wait for Clk_period;
Addr <= "1100101011111";
Trees_din <= "00000000010001010110011000101001";
wait for Clk_period;
Addr <= "1100101100000";
Trees_din <= "00000000001100110110011000101001";
wait for Clk_period;
Addr <= "1100101100001";
Trees_din <= "00000101000000000011101100000100";
wait for Clk_period;
Addr <= "1100101100010";
Trees_din <= "00000000000101000110011000101001";
wait for Clk_period;
Addr <= "1100101100011";
Trees_din <= "00000000010101010110011000101001";
wait for Clk_period;
Addr <= "1100101100100";
Trees_din <= "00000100000000000010000100001000";
wait for Clk_period;
Addr <= "1100101100101";
Trees_din <= "00000110000000000101100000000100";
wait for Clk_period;
Addr <= "1100101100110";
Trees_din <= "00000000010011110110011000101001";
wait for Clk_period;
Addr <= "1100101100111";
Trees_din <= "00000000001001010110011000101001";
wait for Clk_period;
Addr <= "1100101101000";
Trees_din <= "00000110000000000010111000000100";
wait for Clk_period;
Addr <= "1100101101001";
Trees_din <= "00000000000110010110011000101001";
wait for Clk_period;
Addr <= "1100101101010";
Trees_din <= "00000000001001100110011000101001";
wait for Clk_period;
Addr <= "1100101101011";
Trees_din <= "00000101000000000010110100100000";
wait for Clk_period;
Addr <= "1100101101100";
Trees_din <= "00000110000000000001101000010000";
wait for Clk_period;
Addr <= "1100101101101";
Trees_din <= "00000101000000000100011100001000";
wait for Clk_period;
Addr <= "1100101101110";
Trees_din <= "00000010000000000000000100000100";
wait for Clk_period;
Addr <= "1100101101111";
Trees_din <= "00000000010111100110011000101001";
wait for Clk_period;
Addr <= "1100101110000";
Trees_din <= "00000000000111010110011000101001";
wait for Clk_period;
Addr <= "1100101110001";
Trees_din <= "00000001000000000001001000000100";
wait for Clk_period;
Addr <= "1100101110010";
Trees_din <= "00000000001010000110011000101001";
wait for Clk_period;
Addr <= "1100101110011";
Trees_din <= "00000000000000110110011000101001";
wait for Clk_period;
Addr <= "1100101110100";
Trees_din <= "00000110000000000100011100001000";
wait for Clk_period;
Addr <= "1100101110101";
Trees_din <= "00000000000000000011000100000100";
wait for Clk_period;
Addr <= "1100101110110";
Trees_din <= "00000000000001010110011000101001";
wait for Clk_period;
Addr <= "1100101110111";
Trees_din <= "00000000001100100110011000101001";
wait for Clk_period;
Addr <= "1100101111000";
Trees_din <= "00000100000000000100101000000100";
wait for Clk_period;
Addr <= "1100101111001";
Trees_din <= "00000000001100110110011000101001";
wait for Clk_period;
Addr <= "1100101111010";
Trees_din <= "00000000001100000110011000101001";
wait for Clk_period;
Addr <= "1100101111011";
Trees_din <= "00000110000000000001110000010000";
wait for Clk_period;
Addr <= "1100101111100";
Trees_din <= "00000001000000000000110100001000";
wait for Clk_period;
Addr <= "1100101111101";
Trees_din <= "00000111000000000010011000000100";
wait for Clk_period;
Addr <= "1100101111110";
Trees_din <= "00000000000011110110011000101001";
wait for Clk_period;
Addr <= "1100101111111";
Trees_din <= "00000000000000000110011000101001";
wait for Clk_period;
Addr <= "1100110000000";
Trees_din <= "00000100000000000010001100000100";
wait for Clk_period;
Addr <= "1100110000001";
Trees_din <= "00000000001101010110011000101001";
wait for Clk_period;
Addr <= "1100110000010";
Trees_din <= "00000000001111010110011000101001";
wait for Clk_period;
Addr <= "1100110000011";
Trees_din <= "00000010000000000011000100001000";
wait for Clk_period;
Addr <= "1100110000100";
Trees_din <= "00000010000000000100100000000100";
wait for Clk_period;
Addr <= "1100110000101";
Trees_din <= "00000000001100010110011000101001";
wait for Clk_period;
Addr <= "1100110000110";
Trees_din <= "00000000010110110110011000101001";
wait for Clk_period;
Addr <= "1100110000111";
Trees_din <= "00000001000000000100101000000100";
wait for Clk_period;
Addr <= "1100110001000";
Trees_din <= "00000000001100100110011000101001";
wait for Clk_period;
Addr <= "1100110001001";
Trees_din <= "00000000000110000110011000101001";
wait for Clk_period;



----------tree 51-------------------

Addr <= "1100110001010";
Trees_din <= "00000001000000000000001010000000";
wait for Clk_period;
Addr <= "1100110001011";
Trees_din <= "00000110000000000001100001000000";
wait for Clk_period;
Addr <= "1100110001100";
Trees_din <= "00000111000000000100111000100000";
wait for Clk_period;
Addr <= "1100110001101";
Trees_din <= "00000000000000000010101100010000";
wait for Clk_period;
Addr <= "1100110001110";
Trees_din <= "00000011000000000000111000001000";
wait for Clk_period;
Addr <= "1100110001111";
Trees_din <= "00000010000000000001011100000100";
wait for Clk_period;
Addr <= "1100110010000";
Trees_din <= "00000000010100010110100000100101";
wait for Clk_period;
Addr <= "1100110010001";
Trees_din <= "00000000010100100110100000100101";
wait for Clk_period;
Addr <= "1100110010010";
Trees_din <= "00000000000000000011011100000100";
wait for Clk_period;
Addr <= "1100110010011";
Trees_din <= "00000000001000110110100000100101";
wait for Clk_period;
Addr <= "1100110010100";
Trees_din <= "00000000010000100110100000100101";
wait for Clk_period;
Addr <= "1100110010101";
Trees_din <= "00000010000000000000010000001000";
wait for Clk_period;
Addr <= "1100110010110";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "1100110010111";
Trees_din <= "00000000001100000110100000100101";
wait for Clk_period;
Addr <= "1100110011000";
Trees_din <= "00000000000111010110100000100101";
wait for Clk_period;
Addr <= "1100110011001";
Trees_din <= "00000101000000000010000100000100";
wait for Clk_period;
Addr <= "1100110011010";
Trees_din <= "00000000010001010110100000100101";
wait for Clk_period;
Addr <= "1100110011011";
Trees_din <= "00000000000110110110100000100101";
wait for Clk_period;
Addr <= "1100110011100";
Trees_din <= "00000010000000000000000000010000";
wait for Clk_period;
Addr <= "1100110011101";
Trees_din <= "00000001000000000101010000001000";
wait for Clk_period;
Addr <= "1100110011110";
Trees_din <= "00000010000000000100001000000100";
wait for Clk_period;
Addr <= "1100110011111";
Trees_din <= "00000000000111000110100000100101";
wait for Clk_period;
Addr <= "1100110100000";
Trees_din <= "00000000010110100110100000100101";
wait for Clk_period;
Addr <= "1100110100001";
Trees_din <= "00000101000000000000110000000100";
wait for Clk_period;
Addr <= "1100110100010";
Trees_din <= "00000000000011000110100000100101";
wait for Clk_period;
Addr <= "1100110100011";
Trees_din <= "00000000000110000110100000100101";
wait for Clk_period;
Addr <= "1100110100100";
Trees_din <= "00000001000000000101011000001000";
wait for Clk_period;
Addr <= "1100110100101";
Trees_din <= "00000001000000000000011000000100";
wait for Clk_period;
Addr <= "1100110100110";
Trees_din <= "00000000010011110110100000100101";
wait for Clk_period;
Addr <= "1100110100111";
Trees_din <= "00000000001100000110100000100101";
wait for Clk_period;
Addr <= "1100110101000";
Trees_din <= "00000101000000000010101000000100";
wait for Clk_period;
Addr <= "1100110101001";
Trees_din <= "00000000010001110110100000100101";
wait for Clk_period;
Addr <= "1100110101010";
Trees_din <= "00000000000001000110100000100101";
wait for Clk_period;
Addr <= "1100110101011";
Trees_din <= "00000000000000000101000000100000";
wait for Clk_period;
Addr <= "1100110101100";
Trees_din <= "00000001000000000101100000010000";
wait for Clk_period;
Addr <= "1100110101101";
Trees_din <= "00000101000000000100011000001000";
wait for Clk_period;
Addr <= "1100110101110";
Trees_din <= "00000101000000000000011100000100";
wait for Clk_period;
Addr <= "1100110101111";
Trees_din <= "00000000010001000110100000100101";
wait for Clk_period;
Addr <= "1100110110000";
Trees_din <= "00000000000000000110100000100101";
wait for Clk_period;
Addr <= "1100110110001";
Trees_din <= "00000101000000000001111100000100";
wait for Clk_period;
Addr <= "1100110110010";
Trees_din <= "00000000001001110110100000100101";
wait for Clk_period;
Addr <= "1100110110011";
Trees_din <= "00000000010011100110100000100101";
wait for Clk_period;
Addr <= "1100110110100";
Trees_din <= "00000001000000000100100100001000";
wait for Clk_period;
Addr <= "1100110110101";
Trees_din <= "00000011000000000101010100000100";
wait for Clk_period;
Addr <= "1100110110110";
Trees_din <= "00000000010111000110100000100101";
wait for Clk_period;
Addr <= "1100110110111";
Trees_din <= "00000000001110000110100000100101";
wait for Clk_period;
Addr <= "1100110111000";
Trees_din <= "00000111000000000100000000000100";
wait for Clk_period;
Addr <= "1100110111001";
Trees_din <= "00000000001001100110100000100101";
wait for Clk_period;
Addr <= "1100110111010";
Trees_din <= "00000000000011010110100000100101";
wait for Clk_period;
Addr <= "1100110111011";
Trees_din <= "00000100000000000010110100010000";
wait for Clk_period;
Addr <= "1100110111100";
Trees_din <= "00000100000000000011011000001000";
wait for Clk_period;
Addr <= "1100110111101";
Trees_din <= "00000001000000000000101000000100";
wait for Clk_period;
Addr <= "1100110111110";
Trees_din <= "00000000000110110110100000100101";
wait for Clk_period;
Addr <= "1100110111111";
Trees_din <= "00000000010101010110100000100101";
wait for Clk_period;
Addr <= "1100111000000";
Trees_din <= "00000100000000000010000000000100";
wait for Clk_period;
Addr <= "1100111000001";
Trees_din <= "00000000010000010110100000100101";
wait for Clk_period;
Addr <= "1100111000010";
Trees_din <= "00000000011000010110100000100101";
wait for Clk_period;
Addr <= "1100111000011";
Trees_din <= "00000010000000000101010000001000";
wait for Clk_period;
Addr <= "1100111000100";
Trees_din <= "00000000000000000100010100000100";
wait for Clk_period;
Addr <= "1100111000101";
Trees_din <= "00000000010011110110100000100101";
wait for Clk_period;
Addr <= "1100111000110";
Trees_din <= "00000000000010100110100000100101";
wait for Clk_period;
Addr <= "1100111000111";
Trees_din <= "00000101000000000100011100000100";
wait for Clk_period;
Addr <= "1100111001000";
Trees_din <= "00000000001010010110100000100101";
wait for Clk_period;
Addr <= "1100111001001";
Trees_din <= "00000000011001000110100000100101";
wait for Clk_period;
Addr <= "1100111001010";
Trees_din <= "00000010000000000000110101000000";
wait for Clk_period;
Addr <= "1100111001011";
Trees_din <= "00000101000000000100000000100000";
wait for Clk_period;
Addr <= "1100111001100";
Trees_din <= "00000111000000000000110000010000";
wait for Clk_period;
Addr <= "1100111001101";
Trees_din <= "00000010000000000010000000001000";
wait for Clk_period;
Addr <= "1100111001110";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "1100111001111";
Trees_din <= "00000000010101010110100000100101";
wait for Clk_period;
Addr <= "1100111010000";
Trees_din <= "00000000010101000110100000100101";
wait for Clk_period;
Addr <= "1100111010001";
Trees_din <= "00000110000000000010110100000100";
wait for Clk_period;
Addr <= "1100111010010";
Trees_din <= "00000000001000100110100000100101";
wait for Clk_period;
Addr <= "1100111010011";
Trees_din <= "00000000000111000110100000100101";
wait for Clk_period;
Addr <= "1100111010100";
Trees_din <= "00000101000000000101000000001000";
wait for Clk_period;
Addr <= "1100111010101";
Trees_din <= "00000100000000000011000000000100";
wait for Clk_period;
Addr <= "1100111010110";
Trees_din <= "00000000000001110110100000100101";
wait for Clk_period;
Addr <= "1100111010111";
Trees_din <= "00000000001101100110100000100101";
wait for Clk_period;
Addr <= "1100111011000";
Trees_din <= "00000010000000000101001000000100";
wait for Clk_period;
Addr <= "1100111011001";
Trees_din <= "00000000000010110110100000100101";
wait for Clk_period;
Addr <= "1100111011010";
Trees_din <= "00000000000100100110100000100101";
wait for Clk_period;
Addr <= "1100111011011";
Trees_din <= "00000001000000000001010000010000";
wait for Clk_period;
Addr <= "1100111011100";
Trees_din <= "00000011000000000011000100001000";
wait for Clk_period;
Addr <= "1100111011101";
Trees_din <= "00000000000000000110001000000100";
wait for Clk_period;
Addr <= "1100111011110";
Trees_din <= "00000000000111000110100000100101";
wait for Clk_period;
Addr <= "1100111011111";
Trees_din <= "00000000000001100110100000100101";
wait for Clk_period;
Addr <= "1100111100000";
Trees_din <= "00000100000000000101010000000100";
wait for Clk_period;
Addr <= "1100111100001";
Trees_din <= "00000000010010100110100000100101";
wait for Clk_period;
Addr <= "1100111100010";
Trees_din <= "00000000001001000110100000100101";
wait for Clk_period;
Addr <= "1100111100011";
Trees_din <= "00000100000000000101110000001000";
wait for Clk_period;
Addr <= "1100111100100";
Trees_din <= "00000110000000000100100000000100";
wait for Clk_period;
Addr <= "1100111100101";
Trees_din <= "00000000010010110110100000100101";
wait for Clk_period;
Addr <= "1100111100110";
Trees_din <= "00000000010100010110100000100101";
wait for Clk_period;
Addr <= "1100111100111";
Trees_din <= "00000000000000000010001000000100";
wait for Clk_period;
Addr <= "1100111101000";
Trees_din <= "00000000001100010110100000100101";
wait for Clk_period;
Addr <= "1100111101001";
Trees_din <= "00000000001111110110100000100101";
wait for Clk_period;
Addr <= "1100111101010";
Trees_din <= "00000010000000000001001000100000";
wait for Clk_period;
Addr <= "1100111101011";
Trees_din <= "00000111000000000011000100010000";
wait for Clk_period;
Addr <= "1100111101100";
Trees_din <= "00000111000000000000000000001000";
wait for Clk_period;
Addr <= "1100111101101";
Trees_din <= "00000001000000000011010100000100";
wait for Clk_period;
Addr <= "1100111101110";
Trees_din <= "00000000010101110110100000100101";
wait for Clk_period;
Addr <= "1100111101111";
Trees_din <= "00000000011000010110100000100101";
wait for Clk_period;
Addr <= "1100111110000";
Trees_din <= "00000110000000000110000100000100";
wait for Clk_period;
Addr <= "1100111110001";
Trees_din <= "00000000010000010110100000100101";
wait for Clk_period;
Addr <= "1100111110010";
Trees_din <= "00000000010101110110100000100101";
wait for Clk_period;
Addr <= "1100111110011";
Trees_din <= "00000101000000000011010000001000";
wait for Clk_period;
Addr <= "1100111110100";
Trees_din <= "00000111000000000001101000000100";
wait for Clk_period;
Addr <= "1100111110101";
Trees_din <= "00000000000101000110100000100101";
wait for Clk_period;
Addr <= "1100111110110";
Trees_din <= "00000000000111010110100000100101";
wait for Clk_period;
Addr <= "1100111110111";
Trees_din <= "00000111000000000000000000000100";
wait for Clk_period;
Addr <= "1100111111000";
Trees_din <= "00000000010101010110100000100101";
wait for Clk_period;
Addr <= "1100111111001";
Trees_din <= "00000000000100100110100000100101";
wait for Clk_period;
Addr <= "1100111111010";
Trees_din <= "00000000000000000101111100010000";
wait for Clk_period;
Addr <= "1100111111011";
Trees_din <= "00000100000000000100010100001000";
wait for Clk_period;
Addr <= "1100111111100";
Trees_din <= "00000111000000000010010000000100";
wait for Clk_period;
Addr <= "1100111111101";
Trees_din <= "00000000010000100110100000100101";
wait for Clk_period;
Addr <= "1100111111110";
Trees_din <= "00000000000111010110100000100101";
wait for Clk_period;
Addr <= "1100111111111";
Trees_din <= "00000000000000000010111100000100";
wait for Clk_period;
Addr <= "1101000000000";
Trees_din <= "00000000000001110110100000100101";
wait for Clk_period;
Addr <= "1101000000001";
Trees_din <= "00000000010110010110100000100101";
wait for Clk_period;
Addr <= "1101000000010";
Trees_din <= "00000111000000000010000000001000";
wait for Clk_period;
Addr <= "1101000000011";
Trees_din <= "00000001000000000110001100000100";
wait for Clk_period;
Addr <= "1101000000100";
Trees_din <= "00000000001000010110100000100101";
wait for Clk_period;
Addr <= "1101000000101";
Trees_din <= "00000000010000110110100000100101";
wait for Clk_period;
Addr <= "1101000000110";
Trees_din <= "00000000000000000011100100000100";
wait for Clk_period;
Addr <= "1101000000111";
Trees_din <= "00000000010101100110100000100101";
wait for Clk_period;
Addr <= "1101000001000";
Trees_din <= "00000000001001110110100000100101";
wait for Clk_period;



----------tree 52-------------------

Addr <= "1101000001001";
Trees_din <= "00000101000000000100101110000000";
wait for Clk_period;
Addr <= "1101000001010";
Trees_din <= "00000100000000000110010001000000";
wait for Clk_period;
Addr <= "1101000001011";
Trees_din <= "00000100000000000100100000100000";
wait for Clk_period;
Addr <= "1101000001100";
Trees_din <= "00000101000000000011110000010000";
wait for Clk_period;
Addr <= "1101000001101";
Trees_din <= "00000110000000000100100100001000";
wait for Clk_period;
Addr <= "1101000001110";
Trees_din <= "00000010000000000000001100000100";
wait for Clk_period;
Addr <= "1101000001111";
Trees_din <= "00000000001001100110101000100001";
wait for Clk_period;
Addr <= "1101000010000";
Trees_din <= "00000000001001000110101000100001";
wait for Clk_period;
Addr <= "1101000010001";
Trees_din <= "00000000000000000100101000000100";
wait for Clk_period;
Addr <= "1101000010010";
Trees_din <= "00000000011000110110101000100001";
wait for Clk_period;
Addr <= "1101000010011";
Trees_din <= "00000000011000010110101000100001";
wait for Clk_period;
Addr <= "1101000010100";
Trees_din <= "00000010000000000100000000001000";
wait for Clk_period;
Addr <= "1101000010101";
Trees_din <= "00000101000000000100011100000100";
wait for Clk_period;
Addr <= "1101000010110";
Trees_din <= "00000000000100100110101000100001";
wait for Clk_period;
Addr <= "1101000010111";
Trees_din <= "00000000000111010110101000100001";
wait for Clk_period;
Addr <= "1101000011000";
Trees_din <= "00000001000000000011101000000100";
wait for Clk_period;
Addr <= "1101000011001";
Trees_din <= "00000000001011010110101000100001";
wait for Clk_period;
Addr <= "1101000011010";
Trees_din <= "00000000000100010110101000100001";
wait for Clk_period;
Addr <= "1101000011011";
Trees_din <= "00000100000000000100010100010000";
wait for Clk_period;
Addr <= "1101000011100";
Trees_din <= "00000110000000000101100100001000";
wait for Clk_period;
Addr <= "1101000011101";
Trees_din <= "00000011000000000011011000000100";
wait for Clk_period;
Addr <= "1101000011110";
Trees_din <= "00000000001011110110101000100001";
wait for Clk_period;
Addr <= "1101000011111";
Trees_din <= "00000000000110000110101000100001";
wait for Clk_period;
Addr <= "1101000100000";
Trees_din <= "00000010000000000010101000000100";
wait for Clk_period;
Addr <= "1101000100001";
Trees_din <= "00000000011000000110101000100001";
wait for Clk_period;
Addr <= "1101000100010";
Trees_din <= "00000000000110110110101000100001";
wait for Clk_period;
Addr <= "1101000100011";
Trees_din <= "00000011000000000100110000001000";
wait for Clk_period;
Addr <= "1101000100100";
Trees_din <= "00000111000000000100010100000100";
wait for Clk_period;
Addr <= "1101000100101";
Trees_din <= "00000000010010110110101000100001";
wait for Clk_period;
Addr <= "1101000100110";
Trees_din <= "00000000001111010110101000100001";
wait for Clk_period;
Addr <= "1101000100111";
Trees_din <= "00000010000000000101110100000100";
wait for Clk_period;
Addr <= "1101000101000";
Trees_din <= "00000000000000100110101000100001";
wait for Clk_period;
Addr <= "1101000101001";
Trees_din <= "00000000000100000110101000100001";
wait for Clk_period;
Addr <= "1101000101010";
Trees_din <= "00000110000000000010010000100000";
wait for Clk_period;
Addr <= "1101000101011";
Trees_din <= "00000001000000000000010100010000";
wait for Clk_period;
Addr <= "1101000101100";
Trees_din <= "00000011000000000000001000001000";
wait for Clk_period;
Addr <= "1101000101101";
Trees_din <= "00000001000000000000101000000100";
wait for Clk_period;
Addr <= "1101000101110";
Trees_din <= "00000000010110010110101000100001";
wait for Clk_period;
Addr <= "1101000101111";
Trees_din <= "00000000010000000110101000100001";
wait for Clk_period;
Addr <= "1101000110000";
Trees_din <= "00000011000000000100100000000100";
wait for Clk_period;
Addr <= "1101000110001";
Trees_din <= "00000000000111000110101000100001";
wait for Clk_period;
Addr <= "1101000110010";
Trees_din <= "00000000010110010110101000100001";
wait for Clk_period;
Addr <= "1101000110011";
Trees_din <= "00000110000000000001000100001000";
wait for Clk_period;
Addr <= "1101000110100";
Trees_din <= "00000101000000000011111100000100";
wait for Clk_period;
Addr <= "1101000110101";
Trees_din <= "00000000000011010110101000100001";
wait for Clk_period;
Addr <= "1101000110110";
Trees_din <= "00000000001000100110101000100001";
wait for Clk_period;
Addr <= "1101000110111";
Trees_din <= "00000011000000000011110000000100";
wait for Clk_period;
Addr <= "1101000111000";
Trees_din <= "00000000010011010110101000100001";
wait for Clk_period;
Addr <= "1101000111001";
Trees_din <= "00000000000001010110101000100001";
wait for Clk_period;
Addr <= "1101000111010";
Trees_din <= "00000100000000000100111000010000";
wait for Clk_period;
Addr <= "1101000111011";
Trees_din <= "00000011000000000000110100001000";
wait for Clk_period;
Addr <= "1101000111100";
Trees_din <= "00000100000000000010001000000100";
wait for Clk_period;
Addr <= "1101000111101";
Trees_din <= "00000000000000100110101000100001";
wait for Clk_period;
Addr <= "1101000111110";
Trees_din <= "00000000011000010110101000100001";
wait for Clk_period;
Addr <= "1101000111111";
Trees_din <= "00000010000000000101101000000100";
wait for Clk_period;
Addr <= "1101001000000";
Trees_din <= "00000000010101100110101000100001";
wait for Clk_period;
Addr <= "1101001000001";
Trees_din <= "00000000000001100110101000100001";
wait for Clk_period;
Addr <= "1101001000010";
Trees_din <= "00000110000000000011111100001000";
wait for Clk_period;
Addr <= "1101001000011";
Trees_din <= "00000010000000000011110000000100";
wait for Clk_period;
Addr <= "1101001000100";
Trees_din <= "00000000000010010110101000100001";
wait for Clk_period;
Addr <= "1101001000101";
Trees_din <= "00000000001000110110101000100001";
wait for Clk_period;
Addr <= "1101001000110";
Trees_din <= "00000010000000000010100000000100";
wait for Clk_period;
Addr <= "1101001000111";
Trees_din <= "00000000001101000110101000100001";
wait for Clk_period;
Addr <= "1101001001000";
Trees_din <= "00000000000111010110101000100001";
wait for Clk_period;
Addr <= "1101001001001";
Trees_din <= "00000111000000000010101001000000";
wait for Clk_period;
Addr <= "1101001001010";
Trees_din <= "00000011000000000010001100100000";
wait for Clk_period;
Addr <= "1101001001011";
Trees_din <= "00000101000000000100100100010000";
wait for Clk_period;
Addr <= "1101001001100";
Trees_din <= "00000100000000000101101000001000";
wait for Clk_period;
Addr <= "1101001001101";
Trees_din <= "00000010000000000101000000000100";
wait for Clk_period;
Addr <= "1101001001110";
Trees_din <= "00000000011000000110101000100001";
wait for Clk_period;
Addr <= "1101001001111";
Trees_din <= "00000000001111010110101000100001";
wait for Clk_period;
Addr <= "1101001010000";
Trees_din <= "00000010000000000000001000000100";
wait for Clk_period;
Addr <= "1101001010001";
Trees_din <= "00000000010011000110101000100001";
wait for Clk_period;
Addr <= "1101001010010";
Trees_din <= "00000000010000010110101000100001";
wait for Clk_period;
Addr <= "1101001010011";
Trees_din <= "00000011000000000010001000001000";
wait for Clk_period;
Addr <= "1101001010100";
Trees_din <= "00000110000000000011100000000100";
wait for Clk_period;
Addr <= "1101001010101";
Trees_din <= "00000000000101000110101000100001";
wait for Clk_period;
Addr <= "1101001010110";
Trees_din <= "00000000011000000110101000100001";
wait for Clk_period;
Addr <= "1101001010111";
Trees_din <= "00000100000000000100001100000100";
wait for Clk_period;
Addr <= "1101001011000";
Trees_din <= "00000000000100000110101000100001";
wait for Clk_period;
Addr <= "1101001011001";
Trees_din <= "00000000000010100110101000100001";
wait for Clk_period;
Addr <= "1101001011010";
Trees_din <= "00000011000000000110000000010000";
wait for Clk_period;
Addr <= "1101001011011";
Trees_din <= "00000010000000000100010000001000";
wait for Clk_period;
Addr <= "1101001011100";
Trees_din <= "00000110000000000010100100000100";
wait for Clk_period;
Addr <= "1101001011101";
Trees_din <= "00000000000110000110101000100001";
wait for Clk_period;
Addr <= "1101001011110";
Trees_din <= "00000000010010000110101000100001";
wait for Clk_period;
Addr <= "1101001011111";
Trees_din <= "00000111000000000011101100000100";
wait for Clk_period;
Addr <= "1101001100000";
Trees_din <= "00000000000100110110101000100001";
wait for Clk_period;
Addr <= "1101001100001";
Trees_din <= "00000000000010000110101000100001";
wait for Clk_period;
Addr <= "1101001100010";
Trees_din <= "00000100000000000001101000001000";
wait for Clk_period;
Addr <= "1101001100011";
Trees_din <= "00000100000000000010111000000100";
wait for Clk_period;
Addr <= "1101001100100";
Trees_din <= "00000000001000000110101000100001";
wait for Clk_period;
Addr <= "1101001100101";
Trees_din <= "00000000001011010110101000100001";
wait for Clk_period;
Addr <= "1101001100110";
Trees_din <= "00000010000000000100010000000100";
wait for Clk_period;
Addr <= "1101001100111";
Trees_din <= "00000000001001010110101000100001";
wait for Clk_period;
Addr <= "1101001101000";
Trees_din <= "00000000000000100110101000100001";
wait for Clk_period;
Addr <= "1101001101001";
Trees_din <= "00000100000000000001011000100000";
wait for Clk_period;
Addr <= "1101001101010";
Trees_din <= "00000101000000000101100000010000";
wait for Clk_period;
Addr <= "1101001101011";
Trees_din <= "00000111000000000011110100001000";
wait for Clk_period;
Addr <= "1101001101100";
Trees_din <= "00000011000000000011000000000100";
wait for Clk_period;
Addr <= "1101001101101";
Trees_din <= "00000000010010100110101000100001";
wait for Clk_period;
Addr <= "1101001101110";
Trees_din <= "00000000000110000110101000100001";
wait for Clk_period;
Addr <= "1101001101111";
Trees_din <= "00000011000000000110010000000100";
wait for Clk_period;
Addr <= "1101001110000";
Trees_din <= "00000000001110110110101000100001";
wait for Clk_period;
Addr <= "1101001110001";
Trees_din <= "00000000001110010110101000100001";
wait for Clk_period;
Addr <= "1101001110010";
Trees_din <= "00000000000000000000001100001000";
wait for Clk_period;
Addr <= "1101001110011";
Trees_din <= "00000001000000000001100000000100";
wait for Clk_period;
Addr <= "1101001110100";
Trees_din <= "00000000011000010110101000100001";
wait for Clk_period;
Addr <= "1101001110101";
Trees_din <= "00000000001011010110101000100001";
wait for Clk_period;
Addr <= "1101001110110";
Trees_din <= "00000110000000000110001000000100";
wait for Clk_period;
Addr <= "1101001110111";
Trees_din <= "00000000001010110110101000100001";
wait for Clk_period;
Addr <= "1101001111000";
Trees_din <= "00000000010000000110101000100001";
wait for Clk_period;
Addr <= "1101001111001";
Trees_din <= "00000101000000000100001000010000";
wait for Clk_period;
Addr <= "1101001111010";
Trees_din <= "00000110000000000000110000001000";
wait for Clk_period;
Addr <= "1101001111011";
Trees_din <= "00000010000000000010011000000100";
wait for Clk_period;
Addr <= "1101001111100";
Trees_din <= "00000000000001110110101000100001";
wait for Clk_period;
Addr <= "1101001111101";
Trees_din <= "00000000010100000110101000100001";
wait for Clk_period;
Addr <= "1101001111110";
Trees_din <= "00000100000000000000001000000100";
wait for Clk_period;
Addr <= "1101001111111";
Trees_din <= "00000000010001010110101000100001";
wait for Clk_period;
Addr <= "1101010000000";
Trees_din <= "00000000010001000110101000100001";
wait for Clk_period;
Addr <= "1101010000001";
Trees_din <= "00000010000000000101000100001000";
wait for Clk_period;
Addr <= "1101010000010";
Trees_din <= "00000000000000000011110000000100";
wait for Clk_period;
Addr <= "1101010000011";
Trees_din <= "00000000000100100110101000100001";
wait for Clk_period;
Addr <= "1101010000100";
Trees_din <= "00000000001010110110101000100001";
wait for Clk_period;
Addr <= "1101010000101";
Trees_din <= "00000111000000000100001000000100";
wait for Clk_period;
Addr <= "1101010000110";
Trees_din <= "00000000000111000110101000100001";
wait for Clk_period;
Addr <= "1101010000111";
Trees_din <= "00000000010100000110101000100001";
wait for Clk_period;



----------tree 53-------------------

Addr <= "1101010001000";
Trees_din <= "00000011000000000010101110000000";
wait for Clk_period;
Addr <= "1101010001001";
Trees_din <= "00000100000000000100101001000000";
wait for Clk_period;
Addr <= "1101010001010";
Trees_din <= "00000001000000000000100000100000";
wait for Clk_period;
Addr <= "1101010001011";
Trees_din <= "00000000000000000011101100010000";
wait for Clk_period;
Addr <= "1101010001100";
Trees_din <= "00000010000000000011101000001000";
wait for Clk_period;
Addr <= "1101010001101";
Trees_din <= "00000001000000000100111100000100";
wait for Clk_period;
Addr <= "1101010001110";
Trees_din <= "00000000010001100110110000011101";
wait for Clk_period;
Addr <= "1101010001111";
Trees_din <= "00000000010111000110110000011101";
wait for Clk_period;
Addr <= "1101010010000";
Trees_din <= "00000111000000000000111000000100";
wait for Clk_period;
Addr <= "1101010010001";
Trees_din <= "00000000010001110110110000011101";
wait for Clk_period;
Addr <= "1101010010010";
Trees_din <= "00000000001001110110110000011101";
wait for Clk_period;
Addr <= "1101010010011";
Trees_din <= "00000000000000000010011100001000";
wait for Clk_period;
Addr <= "1101010010100";
Trees_din <= "00000010000000000100000100000100";
wait for Clk_period;
Addr <= "1101010010101";
Trees_din <= "00000000000111110110110000011101";
wait for Clk_period;
Addr <= "1101010010110";
Trees_din <= "00000000000010100110110000011101";
wait for Clk_period;
Addr <= "1101010010111";
Trees_din <= "00000010000000000000101100000100";
wait for Clk_period;
Addr <= "1101010011000";
Trees_din <= "00000000010110100110110000011101";
wait for Clk_period;
Addr <= "1101010011001";
Trees_din <= "00000000001101000110110000011101";
wait for Clk_period;
Addr <= "1101010011010";
Trees_din <= "00000100000000000011110100010000";
wait for Clk_period;
Addr <= "1101010011011";
Trees_din <= "00000110000000000100110100001000";
wait for Clk_period;
Addr <= "1101010011100";
Trees_din <= "00000110000000000000010100000100";
wait for Clk_period;
Addr <= "1101010011101";
Trees_din <= "00000000000001000110110000011101";
wait for Clk_period;
Addr <= "1101010011110";
Trees_din <= "00000000010000100110110000011101";
wait for Clk_period;
Addr <= "1101010011111";
Trees_din <= "00000000000000000001000000000100";
wait for Clk_period;
Addr <= "1101010100000";
Trees_din <= "00000000010011110110110000011101";
wait for Clk_period;
Addr <= "1101010100001";
Trees_din <= "00000000001010000110110000011101";
wait for Clk_period;
Addr <= "1101010100010";
Trees_din <= "00000010000000000101100000001000";
wait for Clk_period;
Addr <= "1101010100011";
Trees_din <= "00000100000000000000111100000100";
wait for Clk_period;
Addr <= "1101010100100";
Trees_din <= "00000000001011000110110000011101";
wait for Clk_period;
Addr <= "1101010100101";
Trees_din <= "00000000011000010110110000011101";
wait for Clk_period;
Addr <= "1101010100110";
Trees_din <= "00000001000000000011000000000100";
wait for Clk_period;
Addr <= "1101010100111";
Trees_din <= "00000000000011100110110000011101";
wait for Clk_period;
Addr <= "1101010101000";
Trees_din <= "00000000001000000110110000011101";
wait for Clk_period;
Addr <= "1101010101001";
Trees_din <= "00000011000000000100111100100000";
wait for Clk_period;
Addr <= "1101010101010";
Trees_din <= "00000100000000000100101100010000";
wait for Clk_period;
Addr <= "1101010101011";
Trees_din <= "00000101000000000101000100001000";
wait for Clk_period;
Addr <= "1101010101100";
Trees_din <= "00000011000000000100000000000100";
wait for Clk_period;
Addr <= "1101010101101";
Trees_din <= "00000000001010110110110000011101";
wait for Clk_period;
Addr <= "1101010101110";
Trees_din <= "00000000000001000110110000011101";
wait for Clk_period;
Addr <= "1101010101111";
Trees_din <= "00000110000000000001110000000100";
wait for Clk_period;
Addr <= "1101010110000";
Trees_din <= "00000000011000010110110000011101";
wait for Clk_period;
Addr <= "1101010110001";
Trees_din <= "00000000010111000110110000011101";
wait for Clk_period;
Addr <= "1101010110010";
Trees_din <= "00000110000000000101101100001000";
wait for Clk_period;
Addr <= "1101010110011";
Trees_din <= "00000010000000000100110100000100";
wait for Clk_period;
Addr <= "1101010110100";
Trees_din <= "00000000010101100110110000011101";
wait for Clk_period;
Addr <= "1101010110101";
Trees_din <= "00000000000100110110110000011101";
wait for Clk_period;
Addr <= "1101010110110";
Trees_din <= "00000001000000000010010000000100";
wait for Clk_period;
Addr <= "1101010110111";
Trees_din <= "00000000010111010110110000011101";
wait for Clk_period;
Addr <= "1101010111000";
Trees_din <= "00000000010110000110110000011101";
wait for Clk_period;
Addr <= "1101010111001";
Trees_din <= "00000001000000000100110000010000";
wait for Clk_period;
Addr <= "1101010111010";
Trees_din <= "00000111000000000110001000001000";
wait for Clk_period;
Addr <= "1101010111011";
Trees_din <= "00000111000000000101001000000100";
wait for Clk_period;
Addr <= "1101010111100";
Trees_din <= "00000000001110110110110000011101";
wait for Clk_period;
Addr <= "1101010111101";
Trees_din <= "00000000011001000110110000011101";
wait for Clk_period;
Addr <= "1101010111110";
Trees_din <= "00000001000000000001101000000100";
wait for Clk_period;
Addr <= "1101010111111";
Trees_din <= "00000000010000100110110000011101";
wait for Clk_period;
Addr <= "1101011000000";
Trees_din <= "00000000001101000110110000011101";
wait for Clk_period;
Addr <= "1101011000001";
Trees_din <= "00000001000000000110001100001000";
wait for Clk_period;
Addr <= "1101011000010";
Trees_din <= "00000011000000000011010000000100";
wait for Clk_period;
Addr <= "1101011000011";
Trees_din <= "00000000000011010110110000011101";
wait for Clk_period;
Addr <= "1101011000100";
Trees_din <= "00000000010011000110110000011101";
wait for Clk_period;
Addr <= "1101011000101";
Trees_din <= "00000110000000000100010100000100";
wait for Clk_period;
Addr <= "1101011000110";
Trees_din <= "00000000010010000110110000011101";
wait for Clk_period;
Addr <= "1101011000111";
Trees_din <= "00000000000010110110110000011101";
wait for Clk_period;
Addr <= "1101011001000";
Trees_din <= "00000101000000000011011001000000";
wait for Clk_period;
Addr <= "1101011001001";
Trees_din <= "00000011000000000101001000100000";
wait for Clk_period;
Addr <= "1101011001010";
Trees_din <= "00000001000000000101101000010000";
wait for Clk_period;
Addr <= "1101011001011";
Trees_din <= "00000101000000000100111100001000";
wait for Clk_period;
Addr <= "1101011001100";
Trees_din <= "00000111000000000001001000000100";
wait for Clk_period;
Addr <= "1101011001101";
Trees_din <= "00000000010101000110110000011101";
wait for Clk_period;
Addr <= "1101011001110";
Trees_din <= "00000000010101000110110000011101";
wait for Clk_period;
Addr <= "1101011001111";
Trees_din <= "00000101000000000010100000000100";
wait for Clk_period;
Addr <= "1101011010000";
Trees_din <= "00000000000001000110110000011101";
wait for Clk_period;
Addr <= "1101011010001";
Trees_din <= "00000000000000000110110000011101";
wait for Clk_period;
Addr <= "1101011010010";
Trees_din <= "00000101000000000011001100001000";
wait for Clk_period;
Addr <= "1101011010011";
Trees_din <= "00000010000000000000111100000100";
wait for Clk_period;
Addr <= "1101011010100";
Trees_din <= "00000000000000010110110000011101";
wait for Clk_period;
Addr <= "1101011010101";
Trees_din <= "00000000000100100110110000011101";
wait for Clk_period;
Addr <= "1101011010110";
Trees_din <= "00000100000000000001011100000100";
wait for Clk_period;
Addr <= "1101011010111";
Trees_din <= "00000000010110100110110000011101";
wait for Clk_period;
Addr <= "1101011011000";
Trees_din <= "00000000001111100110110000011101";
wait for Clk_period;
Addr <= "1101011011001";
Trees_din <= "00000001000000000010100000010000";
wait for Clk_period;
Addr <= "1101011011010";
Trees_din <= "00000010000000000010011000001000";
wait for Clk_period;
Addr <= "1101011011011";
Trees_din <= "00000010000000000011101000000100";
wait for Clk_period;
Addr <= "1101011011100";
Trees_din <= "00000000001111100110110000011101";
wait for Clk_period;
Addr <= "1101011011101";
Trees_din <= "00000000001110110110110000011101";
wait for Clk_period;
Addr <= "1101011011110";
Trees_din <= "00000000000000000001111000000100";
wait for Clk_period;
Addr <= "1101011011111";
Trees_din <= "00000000000110010110110000011101";
wait for Clk_period;
Addr <= "1101011100000";
Trees_din <= "00000000000110110110110000011101";
wait for Clk_period;
Addr <= "1101011100001";
Trees_din <= "00000100000000000101111100001000";
wait for Clk_period;
Addr <= "1101011100010";
Trees_din <= "00000101000000000011110000000100";
wait for Clk_period;
Addr <= "1101011100011";
Trees_din <= "00000000010111010110110000011101";
wait for Clk_period;
Addr <= "1101011100100";
Trees_din <= "00000000001100000110110000011101";
wait for Clk_period;
Addr <= "1101011100101";
Trees_din <= "00000100000000000010111000000100";
wait for Clk_period;
Addr <= "1101011100110";
Trees_din <= "00000000001110010110110000011101";
wait for Clk_period;
Addr <= "1101011100111";
Trees_din <= "00000000010101110110110000011101";
wait for Clk_period;
Addr <= "1101011101000";
Trees_din <= "00000111000000000000101000100000";
wait for Clk_period;
Addr <= "1101011101001";
Trees_din <= "00000111000000000100111100010000";
wait for Clk_period;
Addr <= "1101011101010";
Trees_din <= "00000101000000000000010100001000";
wait for Clk_period;
Addr <= "1101011101011";
Trees_din <= "00000000000000000000010000000100";
wait for Clk_period;
Addr <= "1101011101100";
Trees_din <= "00000000010111110110110000011101";
wait for Clk_period;
Addr <= "1101011101101";
Trees_din <= "00000000001101000110110000011101";
wait for Clk_period;
Addr <= "1101011101110";
Trees_din <= "00000101000000000001001000000100";
wait for Clk_period;
Addr <= "1101011101111";
Trees_din <= "00000000000000010110110000011101";
wait for Clk_period;
Addr <= "1101011110000";
Trees_din <= "00000000001101110110110000011101";
wait for Clk_period;
Addr <= "1101011110001";
Trees_din <= "00000011000000000001101100001000";
wait for Clk_period;
Addr <= "1101011110010";
Trees_din <= "00000010000000000100010000000100";
wait for Clk_period;
Addr <= "1101011110011";
Trees_din <= "00000000000011100110110000011101";
wait for Clk_period;
Addr <= "1101011110100";
Trees_din <= "00000000010110110110110000011101";
wait for Clk_period;
Addr <= "1101011110101";
Trees_din <= "00000110000000000101010100000100";
wait for Clk_period;
Addr <= "1101011110110";
Trees_din <= "00000000010001100110110000011101";
wait for Clk_period;
Addr <= "1101011110111";
Trees_din <= "00000000010010000110110000011101";
wait for Clk_period;
Addr <= "1101011111000";
Trees_din <= "00000110000000000000100100010000";
wait for Clk_period;
Addr <= "1101011111001";
Trees_din <= "00000010000000000000011000001000";
wait for Clk_period;
Addr <= "1101011111010";
Trees_din <= "00000001000000000101101100000100";
wait for Clk_period;
Addr <= "1101011111011";
Trees_din <= "00000000001101010110110000011101";
wait for Clk_period;
Addr <= "1101011111100";
Trees_din <= "00000000001000100110110000011101";
wait for Clk_period;
Addr <= "1101011111101";
Trees_din <= "00000101000000000101100000000100";
wait for Clk_period;
Addr <= "1101011111110";
Trees_din <= "00000000011000000110110000011101";
wait for Clk_period;
Addr <= "1101011111111";
Trees_din <= "00000000001000010110110000011101";
wait for Clk_period;
Addr <= "1101100000000";
Trees_din <= "00000001000000000001111000001000";
wait for Clk_period;
Addr <= "1101100000001";
Trees_din <= "00000101000000000000011000000100";
wait for Clk_period;
Addr <= "1101100000010";
Trees_din <= "00000000010001000110110000011101";
wait for Clk_period;
Addr <= "1101100000011";
Trees_din <= "00000000001011000110110000011101";
wait for Clk_period;
Addr <= "1101100000100";
Trees_din <= "00000110000000000001011000000100";
wait for Clk_period;
Addr <= "1101100000101";
Trees_din <= "00000000000110110110110000011101";
wait for Clk_period;
Addr <= "1101100000110";
Trees_din <= "00000000010010010110110000011101";
wait for Clk_period;



----------tree 54-------------------

Addr <= "1101100000111";
Trees_din <= "00000111000000000001110010000000";
wait for Clk_period;
Addr <= "1101100001000";
Trees_din <= "00000001000000000001100101000000";
wait for Clk_period;
Addr <= "1101100001001";
Trees_din <= "00000000000000000001100100100000";
wait for Clk_period;
Addr <= "1101100001010";
Trees_din <= "00000101000000000000110100010000";
wait for Clk_period;
Addr <= "1101100001011";
Trees_din <= "00000010000000000010000100001000";
wait for Clk_period;
Addr <= "1101100001100";
Trees_din <= "00000000000000000001100000000100";
wait for Clk_period;
Addr <= "1101100001101";
Trees_din <= "00000000001111000110111000011011";
wait for Clk_period;
Addr <= "1101100001110";
Trees_din <= "00000000010000110110111000011011";
wait for Clk_period;
Addr <= "1101100001111";
Trees_din <= "00000100000000000101001000000100";
wait for Clk_period;
Addr <= "1101100010000";
Trees_din <= "00000000010000010110111000011011";
wait for Clk_period;
Addr <= "1101100010001";
Trees_din <= "00000000000000110110111000011011";
wait for Clk_period;
Addr <= "1101100010010";
Trees_din <= "00000010000000000100100100001000";
wait for Clk_period;
Addr <= "1101100010011";
Trees_din <= "00000101000000000000100000000100";
wait for Clk_period;
Addr <= "1101100010100";
Trees_din <= "00000000010110010110111000011011";
wait for Clk_period;
Addr <= "1101100010101";
Trees_din <= "00000000001111010110111000011011";
wait for Clk_period;
Addr <= "1101100010110";
Trees_din <= "00000100000000000001101100000100";
wait for Clk_period;
Addr <= "1101100010111";
Trees_din <= "00000000010001110110111000011011";
wait for Clk_period;
Addr <= "1101100011000";
Trees_din <= "00000000000110110110111000011011";
wait for Clk_period;
Addr <= "1101100011001";
Trees_din <= "00000011000000000000001000010000";
wait for Clk_period;
Addr <= "1101100011010";
Trees_din <= "00000100000000000101111000001000";
wait for Clk_period;
Addr <= "1101100011011";
Trees_din <= "00000101000000000001001000000100";
wait for Clk_period;
Addr <= "1101100011100";
Trees_din <= "00000000000100000110111000011011";
wait for Clk_period;
Addr <= "1101100011101";
Trees_din <= "00000000011000100110111000011011";
wait for Clk_period;
Addr <= "1101100011110";
Trees_din <= "00000001000000000100010000000100";
wait for Clk_period;
Addr <= "1101100011111";
Trees_din <= "00000000001001110110111000011011";
wait for Clk_period;
Addr <= "1101100100000";
Trees_din <= "00000000000000100110111000011011";
wait for Clk_period;
Addr <= "1101100100001";
Trees_din <= "00000100000000000110001000001000";
wait for Clk_period;
Addr <= "1101100100010";
Trees_din <= "00000101000000000001000000000100";
wait for Clk_period;
Addr <= "1101100100011";
Trees_din <= "00000000001110010110111000011011";
wait for Clk_period;
Addr <= "1101100100100";
Trees_din <= "00000000001100110110111000011011";
wait for Clk_period;
Addr <= "1101100100101";
Trees_din <= "00000101000000000101010000000100";
wait for Clk_period;
Addr <= "1101100100110";
Trees_din <= "00000000010110000110111000011011";
wait for Clk_period;
Addr <= "1101100100111";
Trees_din <= "00000000010000100110111000011011";
wait for Clk_period;
Addr <= "1101100101000";
Trees_din <= "00000111000000000001010100100000";
wait for Clk_period;
Addr <= "1101100101001";
Trees_din <= "00000111000000000100101000010000";
wait for Clk_period;
Addr <= "1101100101010";
Trees_din <= "00000111000000000100111100001000";
wait for Clk_period;
Addr <= "1101100101011";
Trees_din <= "00000010000000000010000000000100";
wait for Clk_period;
Addr <= "1101100101100";
Trees_din <= "00000000000110000110111000011011";
wait for Clk_period;
Addr <= "1101100101101";
Trees_din <= "00000000010000010110111000011011";
wait for Clk_period;
Addr <= "1101100101110";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "1101100101111";
Trees_din <= "00000000010011010110111000011011";
wait for Clk_period;
Addr <= "1101100110000";
Trees_din <= "00000000001111000110111000011011";
wait for Clk_period;
Addr <= "1101100110001";
Trees_din <= "00000001000000000110010000001000";
wait for Clk_period;
Addr <= "1101100110010";
Trees_din <= "00000010000000000000011100000100";
wait for Clk_period;
Addr <= "1101100110011";
Trees_din <= "00000000011001000110111000011011";
wait for Clk_period;
Addr <= "1101100110100";
Trees_din <= "00000000001110010110111000011011";
wait for Clk_period;
Addr <= "1101100110101";
Trees_din <= "00000001000000000100100100000100";
wait for Clk_period;
Addr <= "1101100110110";
Trees_din <= "00000000000000110110111000011011";
wait for Clk_period;
Addr <= "1101100110111";
Trees_din <= "00000000011000010110111000011011";
wait for Clk_period;
Addr <= "1101100111000";
Trees_din <= "00000110000000000000011100010000";
wait for Clk_period;
Addr <= "1101100111001";
Trees_din <= "00000110000000000000011100001000";
wait for Clk_period;
Addr <= "1101100111010";
Trees_din <= "00000101000000000110010000000100";
wait for Clk_period;
Addr <= "1101100111011";
Trees_din <= "00000000001101000110111000011011";
wait for Clk_period;
Addr <= "1101100111100";
Trees_din <= "00000000000001100110111000011011";
wait for Clk_period;
Addr <= "1101100111101";
Trees_din <= "00000011000000000011110000000100";
wait for Clk_period;
Addr <= "1101100111110";
Trees_din <= "00000000010011010110111000011011";
wait for Clk_period;
Addr <= "1101100111111";
Trees_din <= "00000000010101010110111000011011";
wait for Clk_period;
Addr <= "1101101000000";
Trees_din <= "00000011000000000011100100001000";
wait for Clk_period;
Addr <= "1101101000001";
Trees_din <= "00000001000000000001010100000100";
wait for Clk_period;
Addr <= "1101101000010";
Trees_din <= "00000000010011000110111000011011";
wait for Clk_period;
Addr <= "1101101000011";
Trees_din <= "00000000010111100110111000011011";
wait for Clk_period;
Addr <= "1101101000100";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "1101101000101";
Trees_din <= "00000000000011010110111000011011";
wait for Clk_period;
Addr <= "1101101000110";
Trees_din <= "00000000010010000110111000011011";
wait for Clk_period;
Addr <= "1101101000111";
Trees_din <= "00000111000000000001100001000000";
wait for Clk_period;
Addr <= "1101101001000";
Trees_din <= "00000001000000000010101100100000";
wait for Clk_period;
Addr <= "1101101001001";
Trees_din <= "00000001000000000101111000010000";
wait for Clk_period;
Addr <= "1101101001010";
Trees_din <= "00000010000000000000111100001000";
wait for Clk_period;
Addr <= "1101101001011";
Trees_din <= "00000001000000000100001100000100";
wait for Clk_period;
Addr <= "1101101001100";
Trees_din <= "00000000000000100110111000011011";
wait for Clk_period;
Addr <= "1101101001101";
Trees_din <= "00000000010001010110111000011011";
wait for Clk_period;
Addr <= "1101101001110";
Trees_din <= "00000001000000000001000100000100";
wait for Clk_period;
Addr <= "1101101001111";
Trees_din <= "00000000000010110110111000011011";
wait for Clk_period;
Addr <= "1101101010000";
Trees_din <= "00000000010011000110111000011011";
wait for Clk_period;
Addr <= "1101101010001";
Trees_din <= "00000010000000000010101000001000";
wait for Clk_period;
Addr <= "1101101010010";
Trees_din <= "00000010000000000101110100000100";
wait for Clk_period;
Addr <= "1101101010011";
Trees_din <= "00000000000010000110111000011011";
wait for Clk_period;
Addr <= "1101101010100";
Trees_din <= "00000000011001000110111000011011";
wait for Clk_period;
Addr <= "1101101010101";
Trees_din <= "00000110000000000101000000000100";
wait for Clk_period;
Addr <= "1101101010110";
Trees_din <= "00000000010011100110111000011011";
wait for Clk_period;
Addr <= "1101101010111";
Trees_din <= "00000000001010000110111000011011";
wait for Clk_period;
Addr <= "1101101011000";
Trees_din <= "00000010000000000010100000010000";
wait for Clk_period;
Addr <= "1101101011001";
Trees_din <= "00000101000000000000000100001000";
wait for Clk_period;
Addr <= "1101101011010";
Trees_din <= "00000001000000000010011000000100";
wait for Clk_period;
Addr <= "1101101011011";
Trees_din <= "00000000000011110110111000011011";
wait for Clk_period;
Addr <= "1101101011100";
Trees_din <= "00000000001001000110111000011011";
wait for Clk_period;
Addr <= "1101101011101";
Trees_din <= "00000100000000000100001100000100";
wait for Clk_period;
Addr <= "1101101011110";
Trees_din <= "00000000011000100110111000011011";
wait for Clk_period;
Addr <= "1101101011111";
Trees_din <= "00000000010100000110111000011011";
wait for Clk_period;
Addr <= "1101101100000";
Trees_din <= "00000111000000000001110000001000";
wait for Clk_period;
Addr <= "1101101100001";
Trees_din <= "00000100000000000101000000000100";
wait for Clk_period;
Addr <= "1101101100010";
Trees_din <= "00000000000001010110111000011011";
wait for Clk_period;
Addr <= "1101101100011";
Trees_din <= "00000000010101110110111000011011";
wait for Clk_period;
Addr <= "1101101100100";
Trees_din <= "00000101000000000000000100000100";
wait for Clk_period;
Addr <= "1101101100101";
Trees_din <= "00000000010011110110111000011011";
wait for Clk_period;
Addr <= "1101101100110";
Trees_din <= "00000000010111000110111000011011";
wait for Clk_period;
Addr <= "1101101100111";
Trees_din <= "00000101000000000101101100100000";
wait for Clk_period;
Addr <= "1101101101000";
Trees_din <= "00000000000000000001011000010000";
wait for Clk_period;
Addr <= "1101101101001";
Trees_din <= "00000000000000000000001100001000";
wait for Clk_period;
Addr <= "1101101101010";
Trees_din <= "00000111000000000011100100000100";
wait for Clk_period;
Addr <= "1101101101011";
Trees_din <= "00000000001100010110111000011011";
wait for Clk_period;
Addr <= "1101101101100";
Trees_din <= "00000000001100100110111000011011";
wait for Clk_period;
Addr <= "1101101101101";
Trees_din <= "00000101000000000001110100000100";
wait for Clk_period;
Addr <= "1101101101110";
Trees_din <= "00000000010111100110111000011011";
wait for Clk_period;
Addr <= "1101101101111";
Trees_din <= "00000000001000110110111000011011";
wait for Clk_period;
Addr <= "1101101110000";
Trees_din <= "00000011000000000100101000001000";
wait for Clk_period;
Addr <= "1101101110001";
Trees_din <= "00000101000000000001011100000100";
wait for Clk_period;
Addr <= "1101101110010";
Trees_din <= "00000000010000110110111000011011";
wait for Clk_period;
Addr <= "1101101110011";
Trees_din <= "00000000001101000110111000011011";
wait for Clk_period;
Addr <= "1101101110100";
Trees_din <= "00000110000000000010010000000100";
wait for Clk_period;
Addr <= "1101101110101";
Trees_din <= "00000000010110000110111000011011";
wait for Clk_period;
Addr <= "1101101110110";
Trees_din <= "00000000001111100110111000011011";
wait for Clk_period;
Addr <= "1101101110111";
Trees_din <= "00000100000000000101111000010000";
wait for Clk_period;
Addr <= "1101101111000";
Trees_din <= "00000000000000000000100000001000";
wait for Clk_period;
Addr <= "1101101111001";
Trees_din <= "00000011000000000000101100000100";
wait for Clk_period;
Addr <= "1101101111010";
Trees_din <= "00000000000011100110111000011011";
wait for Clk_period;
Addr <= "1101101111011";
Trees_din <= "00000000000001100110111000011011";
wait for Clk_period;
Addr <= "1101101111100";
Trees_din <= "00000100000000000011100000000100";
wait for Clk_period;
Addr <= "1101101111101";
Trees_din <= "00000000000010110110111000011011";
wait for Clk_period;
Addr <= "1101101111110";
Trees_din <= "00000000001010100110111000011011";
wait for Clk_period;
Addr <= "1101101111111";
Trees_din <= "00000101000000000101110000001000";
wait for Clk_period;
Addr <= "1101110000000";
Trees_din <= "00000000000000000101010100000100";
wait for Clk_period;
Addr <= "1101110000001";
Trees_din <= "00000000010010110110111000011011";
wait for Clk_period;
Addr <= "1101110000010";
Trees_din <= "00000000001011010110111000011011";
wait for Clk_period;
Addr <= "1101110000011";
Trees_din <= "00000001000000000100000000000100";
wait for Clk_period;
Addr <= "1101110000100";
Trees_din <= "00000000000000100110111000011011";
wait for Clk_period;
Addr <= "1101110000101";
Trees_din <= "00000000000110110110111000011011";
wait for Clk_period;



----------tree 55-------------------

Addr <= "1101110000110";
Trees_din <= "00000100000000000001011010000000";
wait for Clk_period;
Addr <= "1101110000111";
Trees_din <= "00000000000000000100111101000000";
wait for Clk_period;
Addr <= "1101110001000";
Trees_din <= "00000110000000000101001100100000";
wait for Clk_period;
Addr <= "1101110001001";
Trees_din <= "00000001000000000000100000010000";
wait for Clk_period;
Addr <= "1101110001010";
Trees_din <= "00000010000000000100011000001000";
wait for Clk_period;
Addr <= "1101110001011";
Trees_din <= "00000001000000000101100000000100";
wait for Clk_period;
Addr <= "1101110001100";
Trees_din <= "00000000010001010111000000010101";
wait for Clk_period;
Addr <= "1101110001101";
Trees_din <= "00000000000100010111000000010101";
wait for Clk_period;
Addr <= "1101110001110";
Trees_din <= "00000110000000000100010100000100";
wait for Clk_period;
Addr <= "1101110001111";
Trees_din <= "00000000000100010111000000010101";
wait for Clk_period;
Addr <= "1101110010000";
Trees_din <= "00000000010111000111000000010101";
wait for Clk_period;
Addr <= "1101110010001";
Trees_din <= "00000111000000000000000000001000";
wait for Clk_period;
Addr <= "1101110010010";
Trees_din <= "00000110000000000010100100000100";
wait for Clk_period;
Addr <= "1101110010011";
Trees_din <= "00000000011000110111000000010101";
wait for Clk_period;
Addr <= "1101110010100";
Trees_din <= "00000000010010100111000000010101";
wait for Clk_period;
Addr <= "1101110010101";
Trees_din <= "00000011000000000010010100000100";
wait for Clk_period;
Addr <= "1101110010110";
Trees_din <= "00000000001001110111000000010101";
wait for Clk_period;
Addr <= "1101110010111";
Trees_din <= "00000000001110010111000000010101";
wait for Clk_period;
Addr <= "1101110011000";
Trees_din <= "00000001000000000000100100010000";
wait for Clk_period;
Addr <= "1101110011001";
Trees_din <= "00000011000000000110000100001000";
wait for Clk_period;
Addr <= "1101110011010";
Trees_din <= "00000100000000000011011100000100";
wait for Clk_period;
Addr <= "1101110011011";
Trees_din <= "00000000010100100111000000010101";
wait for Clk_period;
Addr <= "1101110011100";
Trees_din <= "00000000001101110111000000010101";
wait for Clk_period;
Addr <= "1101110011101";
Trees_din <= "00000100000000000011000000000100";
wait for Clk_period;
Addr <= "1101110011110";
Trees_din <= "00000000010111100111000000010101";
wait for Clk_period;
Addr <= "1101110011111";
Trees_din <= "00000000010001000111000000010101";
wait for Clk_period;
Addr <= "1101110100000";
Trees_din <= "00000000000000000010111100001000";
wait for Clk_period;
Addr <= "1101110100001";
Trees_din <= "00000100000000000001111000000100";
wait for Clk_period;
Addr <= "1101110100010";
Trees_din <= "00000000000101100111000000010101";
wait for Clk_period;
Addr <= "1101110100011";
Trees_din <= "00000000011000100111000000010101";
wait for Clk_period;
Addr <= "1101110100100";
Trees_din <= "00000100000000000000000000000100";
wait for Clk_period;
Addr <= "1101110100101";
Trees_din <= "00000000001100000111000000010101";
wait for Clk_period;
Addr <= "1101110100110";
Trees_din <= "00000000000101010111000000010101";
wait for Clk_period;
Addr <= "1101110100111";
Trees_din <= "00000000000000000010001100100000";
wait for Clk_period;
Addr <= "1101110101000";
Trees_din <= "00000010000000000000010000010000";
wait for Clk_period;
Addr <= "1101110101001";
Trees_din <= "00000111000000000010111000001000";
wait for Clk_period;
Addr <= "1101110101010";
Trees_din <= "00000010000000000010101100000100";
wait for Clk_period;
Addr <= "1101110101011";
Trees_din <= "00000000010010110111000000010101";
wait for Clk_period;
Addr <= "1101110101100";
Trees_din <= "00000000010000000111000000010101";
wait for Clk_period;
Addr <= "1101110101101";
Trees_din <= "00000110000000000101101100000100";
wait for Clk_period;
Addr <= "1101110101110";
Trees_din <= "00000000001011110111000000010101";
wait for Clk_period;
Addr <= "1101110101111";
Trees_din <= "00000000001101100111000000010101";
wait for Clk_period;
Addr <= "1101110110000";
Trees_din <= "00000001000000000010011000001000";
wait for Clk_period;
Addr <= "1101110110001";
Trees_din <= "00000100000000000000100100000100";
wait for Clk_period;
Addr <= "1101110110010";
Trees_din <= "00000000010011010111000000010101";
wait for Clk_period;
Addr <= "1101110110011";
Trees_din <= "00000000000101000111000000010101";
wait for Clk_period;
Addr <= "1101110110100";
Trees_din <= "00000110000000000100010000000100";
wait for Clk_period;
Addr <= "1101110110101";
Trees_din <= "00000000000010000111000000010101";
wait for Clk_period;
Addr <= "1101110110110";
Trees_din <= "00000000010011010111000000010101";
wait for Clk_period;
Addr <= "1101110110111";
Trees_din <= "00000100000000000000101100010000";
wait for Clk_period;
Addr <= "1101110111000";
Trees_din <= "00000000000000000001111100001000";
wait for Clk_period;
Addr <= "1101110111001";
Trees_din <= "00000010000000000011010000000100";
wait for Clk_period;
Addr <= "1101110111010";
Trees_din <= "00000000010000110111000000010101";
wait for Clk_period;
Addr <= "1101110111011";
Trees_din <= "00000000000101110111000000010101";
wait for Clk_period;
Addr <= "1101110111100";
Trees_din <= "00000000000000000011010000000100";
wait for Clk_period;
Addr <= "1101110111101";
Trees_din <= "00000000000111010111000000010101";
wait for Clk_period;
Addr <= "1101110111110";
Trees_din <= "00000000010000100111000000010101";
wait for Clk_period;
Addr <= "1101110111111";
Trees_din <= "00000100000000000010000100001000";
wait for Clk_period;
Addr <= "1101111000000";
Trees_din <= "00000110000000000100111100000100";
wait for Clk_period;
Addr <= "1101111000001";
Trees_din <= "00000000000111000111000000010101";
wait for Clk_period;
Addr <= "1101111000010";
Trees_din <= "00000000001110010111000000010101";
wait for Clk_period;
Addr <= "1101111000011";
Trees_din <= "00000110000000000011011000000100";
wait for Clk_period;
Addr <= "1101111000100";
Trees_din <= "00000000001000110111000000010101";
wait for Clk_period;
Addr <= "1101111000101";
Trees_din <= "00000000000000100111000000010101";
wait for Clk_period;
Addr <= "1101111000110";
Trees_din <= "00000100000000000100011101000000";
wait for Clk_period;
Addr <= "1101111000111";
Trees_din <= "00000110000000000000100000100000";
wait for Clk_period;
Addr <= "1101111001000";
Trees_din <= "00000100000000000010001100010000";
wait for Clk_period;
Addr <= "1101111001001";
Trees_din <= "00000110000000000011000100001000";
wait for Clk_period;
Addr <= "1101111001010";
Trees_din <= "00000100000000000100111000000100";
wait for Clk_period;
Addr <= "1101111001011";
Trees_din <= "00000000000010010111000000010101";
wait for Clk_period;
Addr <= "1101111001100";
Trees_din <= "00000000000110010111000000010101";
wait for Clk_period;
Addr <= "1101111001101";
Trees_din <= "00000011000000000011001100000100";
wait for Clk_period;
Addr <= "1101111001110";
Trees_din <= "00000000000110000111000000010101";
wait for Clk_period;
Addr <= "1101111001111";
Trees_din <= "00000000000101010111000000010101";
wait for Clk_period;
Addr <= "1101111010000";
Trees_din <= "00000111000000000011110000001000";
wait for Clk_period;
Addr <= "1101111010001";
Trees_din <= "00000101000000000110001000000100";
wait for Clk_period;
Addr <= "1101111010010";
Trees_din <= "00000000001010000111000000010101";
wait for Clk_period;
Addr <= "1101111010011";
Trees_din <= "00000000010100000111000000010101";
wait for Clk_period;
Addr <= "1101111010100";
Trees_din <= "00000010000000000000100100000100";
wait for Clk_period;
Addr <= "1101111010101";
Trees_din <= "00000000000000110111000000010101";
wait for Clk_period;
Addr <= "1101111010110";
Trees_din <= "00000000010010100111000000010101";
wait for Clk_period;
Addr <= "1101111010111";
Trees_din <= "00000111000000000001110100010000";
wait for Clk_period;
Addr <= "1101111011000";
Trees_din <= "00000111000000000001001100001000";
wait for Clk_period;
Addr <= "1101111011001";
Trees_din <= "00000000000000000100110000000100";
wait for Clk_period;
Addr <= "1101111011010";
Trees_din <= "00000000000011010111000000010101";
wait for Clk_period;
Addr <= "1101111011011";
Trees_din <= "00000000000111110111000000010101";
wait for Clk_period;
Addr <= "1101111011100";
Trees_din <= "00000110000000000000110100000100";
wait for Clk_period;
Addr <= "1101111011101";
Trees_din <= "00000000001001000111000000010101";
wait for Clk_period;
Addr <= "1101111011110";
Trees_din <= "00000000000010010111000000010101";
wait for Clk_period;
Addr <= "1101111011111";
Trees_din <= "00000100000000000011100000001000";
wait for Clk_period;
Addr <= "1101111100000";
Trees_din <= "00000101000000000001011100000100";
wait for Clk_period;
Addr <= "1101111100001";
Trees_din <= "00000000010101000111000000010101";
wait for Clk_period;
Addr <= "1101111100010";
Trees_din <= "00000000010110000111000000010101";
wait for Clk_period;
Addr <= "1101111100011";
Trees_din <= "00000111000000000000100100000100";
wait for Clk_period;
Addr <= "1101111100100";
Trees_din <= "00000000011001000111000000010101";
wait for Clk_period;
Addr <= "1101111100101";
Trees_din <= "00000000010000110111000000010101";
wait for Clk_period;
Addr <= "1101111100110";
Trees_din <= "00000010000000000010100000100000";
wait for Clk_period;
Addr <= "1101111100111";
Trees_din <= "00000011000000000110010000010000";
wait for Clk_period;
Addr <= "1101111101000";
Trees_din <= "00000110000000000100000000001000";
wait for Clk_period;
Addr <= "1101111101001";
Trees_din <= "00000101000000000011111000000100";
wait for Clk_period;
Addr <= "1101111101010";
Trees_din <= "00000000010101100111000000010101";
wait for Clk_period;
Addr <= "1101111101011";
Trees_din <= "00000000010111010111000000010101";
wait for Clk_period;
Addr <= "1101111101100";
Trees_din <= "00000101000000000101100100000100";
wait for Clk_period;
Addr <= "1101111101101";
Trees_din <= "00000000001101010111000000010101";
wait for Clk_period;
Addr <= "1101111101110";
Trees_din <= "00000000010010000111000000010101";
wait for Clk_period;
Addr <= "1101111101111";
Trees_din <= "00000101000000000100010100001000";
wait for Clk_period;
Addr <= "1101111110000";
Trees_din <= "00000101000000000000100000000100";
wait for Clk_period;
Addr <= "1101111110001";
Trees_din <= "00000000010011100111000000010101";
wait for Clk_period;
Addr <= "1101111110010";
Trees_din <= "00000000000010010111000000010101";
wait for Clk_period;
Addr <= "1101111110011";
Trees_din <= "00000100000000000000001000000100";
wait for Clk_period;
Addr <= "1101111110100";
Trees_din <= "00000000001010000111000000010101";
wait for Clk_period;
Addr <= "1101111110101";
Trees_din <= "00000000001010000111000000010101";
wait for Clk_period;
Addr <= "1101111110110";
Trees_din <= "00000010000000000101110100010000";
wait for Clk_period;
Addr <= "1101111110111";
Trees_din <= "00000101000000000000110000001000";
wait for Clk_period;
Addr <= "1101111111000";
Trees_din <= "00000111000000000101100000000100";
wait for Clk_period;
Addr <= "1101111111001";
Trees_din <= "00000000000011100111000000010101";
wait for Clk_period;
Addr <= "1101111111010";
Trees_din <= "00000000010110000111000000010101";
wait for Clk_period;
Addr <= "1101111111011";
Trees_din <= "00000000000000000010100100000100";
wait for Clk_period;
Addr <= "1101111111100";
Trees_din <= "00000000000111010111000000010101";
wait for Clk_period;
Addr <= "1101111111101";
Trees_din <= "00000000001010010111000000010101";
wait for Clk_period;
Addr <= "1101111111110";
Trees_din <= "00000101000000000101010100001000";
wait for Clk_period;
Addr <= "1101111111111";
Trees_din <= "00000100000000000100010100000100";
wait for Clk_period;
Addr <= "1110000000000";
Trees_din <= "00000000010010000111000000010101";
wait for Clk_period;
Addr <= "1110000000001";
Trees_din <= "00000000001111000111000000010101";
wait for Clk_period;
Addr <= "1110000000010";
Trees_din <= "00000011000000000100111000000100";
wait for Clk_period;
Addr <= "1110000000011";
Trees_din <= "00000000010011100111000000010101";
wait for Clk_period;
Addr <= "1110000000100";
Trees_din <= "00000000010001010111000000010101";
wait for Clk_period;



----------tree 56-------------------

Addr <= "1110000000101";
Trees_din <= "00000101000000000100011010000000";
wait for Clk_period;
Addr <= "1110000000110";
Trees_din <= "00000101000000000010000101000000";
wait for Clk_period;
Addr <= "1110000000111";
Trees_din <= "00000110000000000000111000100000";
wait for Clk_period;
Addr <= "1110000001000";
Trees_din <= "00000100000000000101101000010000";
wait for Clk_period;
Addr <= "1110000001001";
Trees_din <= "00000001000000000001011000001000";
wait for Clk_period;
Addr <= "1110000001010";
Trees_din <= "00000100000000000101111100000100";
wait for Clk_period;
Addr <= "1110000001011";
Trees_din <= "00000000001110000111001000010001";
wait for Clk_period;
Addr <= "1110000001100";
Trees_din <= "00000000001001000111001000010001";
wait for Clk_period;
Addr <= "1110000001101";
Trees_din <= "00000100000000000100011000000100";
wait for Clk_period;
Addr <= "1110000001110";
Trees_din <= "00000000010000010111001000010001";
wait for Clk_period;
Addr <= "1110000001111";
Trees_din <= "00000000010010010111001000010001";
wait for Clk_period;
Addr <= "1110000010000";
Trees_din <= "00000111000000000000010000001000";
wait for Clk_period;
Addr <= "1110000010001";
Trees_din <= "00000011000000000011100000000100";
wait for Clk_period;
Addr <= "1110000010010";
Trees_din <= "00000000000101000111001000010001";
wait for Clk_period;
Addr <= "1110000010011";
Trees_din <= "00000000010000000111001000010001";
wait for Clk_period;
Addr <= "1110000010100";
Trees_din <= "00000001000000000001110100000100";
wait for Clk_period;
Addr <= "1110000010101";
Trees_din <= "00000000001010010111001000010001";
wait for Clk_period;
Addr <= "1110000010110";
Trees_din <= "00000000000110000111001000010001";
wait for Clk_period;
Addr <= "1110000010111";
Trees_din <= "00000110000000000100110100010000";
wait for Clk_period;
Addr <= "1110000011000";
Trees_din <= "00000000000000000000001000001000";
wait for Clk_period;
Addr <= "1110000011001";
Trees_din <= "00000110000000000101101100000100";
wait for Clk_period;
Addr <= "1110000011010";
Trees_din <= "00000000010101110111001000010001";
wait for Clk_period;
Addr <= "1110000011011";
Trees_din <= "00000000010011100111001000010001";
wait for Clk_period;
Addr <= "1110000011100";
Trees_din <= "00000011000000000001110000000100";
wait for Clk_period;
Addr <= "1110000011101";
Trees_din <= "00000000000011000111001000010001";
wait for Clk_period;
Addr <= "1110000011110";
Trees_din <= "00000000000100000111001000010001";
wait for Clk_period;
Addr <= "1110000011111";
Trees_din <= "00000011000000000100110100001000";
wait for Clk_period;
Addr <= "1110000100000";
Trees_din <= "00000101000000000001111000000100";
wait for Clk_period;
Addr <= "1110000100001";
Trees_din <= "00000000001110100111001000010001";
wait for Clk_period;
Addr <= "1110000100010";
Trees_din <= "00000000001110110111001000010001";
wait for Clk_period;
Addr <= "1110000100011";
Trees_din <= "00000001000000000101111000000100";
wait for Clk_period;
Addr <= "1110000100100";
Trees_din <= "00000000010001110111001000010001";
wait for Clk_period;
Addr <= "1110000100101";
Trees_din <= "00000000000000100111001000010001";
wait for Clk_period;
Addr <= "1110000100110";
Trees_din <= "00000111000000000001101100100000";
wait for Clk_period;
Addr <= "1110000100111";
Trees_din <= "00000001000000000101110100010000";
wait for Clk_period;
Addr <= "1110000101000";
Trees_din <= "00000001000000000000100000001000";
wait for Clk_period;
Addr <= "1110000101001";
Trees_din <= "00000011000000000010101100000100";
wait for Clk_period;
Addr <= "1110000101010";
Trees_din <= "00000000010100110111001000010001";
wait for Clk_period;
Addr <= "1110000101011";
Trees_din <= "00000000001000000111001000010001";
wait for Clk_period;
Addr <= "1110000101100";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "1110000101101";
Trees_din <= "00000000001010100111001000010001";
wait for Clk_period;
Addr <= "1110000101110";
Trees_din <= "00000000010101100111001000010001";
wait for Clk_period;
Addr <= "1110000101111";
Trees_din <= "00000000000000000011110000001000";
wait for Clk_period;
Addr <= "1110000110000";
Trees_din <= "00000111000000000000010000000100";
wait for Clk_period;
Addr <= "1110000110001";
Trees_din <= "00000000001011010111001000010001";
wait for Clk_period;
Addr <= "1110000110010";
Trees_din <= "00000000000101000111001000010001";
wait for Clk_period;
Addr <= "1110000110011";
Trees_din <= "00000010000000000000000000000100";
wait for Clk_period;
Addr <= "1110000110100";
Trees_din <= "00000000000101010111001000010001";
wait for Clk_period;
Addr <= "1110000110101";
Trees_din <= "00000000010110000111001000010001";
wait for Clk_period;
Addr <= "1110000110110";
Trees_din <= "00000001000000000000101100010000";
wait for Clk_period;
Addr <= "1110000110111";
Trees_din <= "00000110000000000000111000001000";
wait for Clk_period;
Addr <= "1110000111000";
Trees_din <= "00000000000000000001010100000100";
wait for Clk_period;
Addr <= "1110000111001";
Trees_din <= "00000000000101000111001000010001";
wait for Clk_period;
Addr <= "1110000111010";
Trees_din <= "00000000000100010111001000010001";
wait for Clk_period;
Addr <= "1110000111011";
Trees_din <= "00000100000000000011101000000100";
wait for Clk_period;
Addr <= "1110000111100";
Trees_din <= "00000000010100110111001000010001";
wait for Clk_period;
Addr <= "1110000111101";
Trees_din <= "00000000010101010111001000010001";
wait for Clk_period;
Addr <= "1110000111110";
Trees_din <= "00000010000000000011001100001000";
wait for Clk_period;
Addr <= "1110000111111";
Trees_din <= "00000110000000000101000000000100";
wait for Clk_period;
Addr <= "1110001000000";
Trees_din <= "00000000010011000111001000010001";
wait for Clk_period;
Addr <= "1110001000001";
Trees_din <= "00000000010110010111001000010001";
wait for Clk_period;
Addr <= "1110001000010";
Trees_din <= "00000011000000000101111000000100";
wait for Clk_period;
Addr <= "1110001000011";
Trees_din <= "00000000010100000111001000010001";
wait for Clk_period;
Addr <= "1110001000100";
Trees_din <= "00000000010101000111001000010001";
wait for Clk_period;
Addr <= "1110001000101";
Trees_din <= "00000001000000000100001001000000";
wait for Clk_period;
Addr <= "1110001000110";
Trees_din <= "00000100000000000100011100100000";
wait for Clk_period;
Addr <= "1110001000111";
Trees_din <= "00000001000000000100011000010000";
wait for Clk_period;
Addr <= "1110001001000";
Trees_din <= "00000001000000000101111000001000";
wait for Clk_period;
Addr <= "1110001001001";
Trees_din <= "00000001000000000101110100000100";
wait for Clk_period;
Addr <= "1110001001010";
Trees_din <= "00000000000101110111001000010001";
wait for Clk_period;
Addr <= "1110001001011";
Trees_din <= "00000000010010110111001000010001";
wait for Clk_period;
Addr <= "1110001001100";
Trees_din <= "00000000000000000110010000000100";
wait for Clk_period;
Addr <= "1110001001101";
Trees_din <= "00000000000101100111001000010001";
wait for Clk_period;
Addr <= "1110001001110";
Trees_din <= "00000000001010100111001000010001";
wait for Clk_period;
Addr <= "1110001001111";
Trees_din <= "00000010000000000000000100001000";
wait for Clk_period;
Addr <= "1110001010000";
Trees_din <= "00000010000000000001101100000100";
wait for Clk_period;
Addr <= "1110001010001";
Trees_din <= "00000000010011110111001000010001";
wait for Clk_period;
Addr <= "1110001010010";
Trees_din <= "00000000010111000111001000010001";
wait for Clk_period;
Addr <= "1110001010011";
Trees_din <= "00000111000000000010011000000100";
wait for Clk_period;
Addr <= "1110001010100";
Trees_din <= "00000000010100100111001000010001";
wait for Clk_period;
Addr <= "1110001010101";
Trees_din <= "00000000001100000111001000010001";
wait for Clk_period;
Addr <= "1110001010110";
Trees_din <= "00000001000000000001110100010000";
wait for Clk_period;
Addr <= "1110001010111";
Trees_din <= "00000011000000000100010100001000";
wait for Clk_period;
Addr <= "1110001011000";
Trees_din <= "00000101000000000010111100000100";
wait for Clk_period;
Addr <= "1110001011001";
Trees_din <= "00000000010001010111001000010001";
wait for Clk_period;
Addr <= "1110001011010";
Trees_din <= "00000000001011100111001000010001";
wait for Clk_period;
Addr <= "1110001011011";
Trees_din <= "00000011000000000001101100000100";
wait for Clk_period;
Addr <= "1110001011100";
Trees_din <= "00000000001101100111001000010001";
wait for Clk_period;
Addr <= "1110001011101";
Trees_din <= "00000000010011100111001000010001";
wait for Clk_period;
Addr <= "1110001011110";
Trees_din <= "00000111000000000101011100001000";
wait for Clk_period;
Addr <= "1110001011111";
Trees_din <= "00000000000000000000010000000100";
wait for Clk_period;
Addr <= "1110001100000";
Trees_din <= "00000000000011110111001000010001";
wait for Clk_period;
Addr <= "1110001100001";
Trees_din <= "00000000000111100111001000010001";
wait for Clk_period;
Addr <= "1110001100010";
Trees_din <= "00000110000000000010100100000100";
wait for Clk_period;
Addr <= "1110001100011";
Trees_din <= "00000000011000010111001000010001";
wait for Clk_period;
Addr <= "1110001100100";
Trees_din <= "00000000001001010111001000010001";
wait for Clk_period;
Addr <= "1110001100101";
Trees_din <= "00000010000000000010001100100000";
wait for Clk_period;
Addr <= "1110001100110";
Trees_din <= "00000101000000000001010000010000";
wait for Clk_period;
Addr <= "1110001100111";
Trees_din <= "00000000000000000010000100001000";
wait for Clk_period;
Addr <= "1110001101000";
Trees_din <= "00000101000000000011010000000100";
wait for Clk_period;
Addr <= "1110001101001";
Trees_din <= "00000000001111010111001000010001";
wait for Clk_period;
Addr <= "1110001101010";
Trees_din <= "00000000000101000111001000010001";
wait for Clk_period;
Addr <= "1110001101011";
Trees_din <= "00000110000000000000111100000100";
wait for Clk_period;
Addr <= "1110001101100";
Trees_din <= "00000000000100110111001000010001";
wait for Clk_period;
Addr <= "1110001101101";
Trees_din <= "00000000010011110111001000010001";
wait for Clk_period;
Addr <= "1110001101110";
Trees_din <= "00000000000000000100000000001000";
wait for Clk_period;
Addr <= "1110001101111";
Trees_din <= "00000000000000000101111000000100";
wait for Clk_period;
Addr <= "1110001110000";
Trees_din <= "00000000010000100111001000010001";
wait for Clk_period;
Addr <= "1110001110001";
Trees_din <= "00000000010110010111001000010001";
wait for Clk_period;
Addr <= "1110001110010";
Trees_din <= "00000101000000000001010000000100";
wait for Clk_period;
Addr <= "1110001110011";
Trees_din <= "00000000010101100111001000010001";
wait for Clk_period;
Addr <= "1110001110100";
Trees_din <= "00000000010011010111001000010001";
wait for Clk_period;
Addr <= "1110001110101";
Trees_din <= "00000010000000000100101000010000";
wait for Clk_period;
Addr <= "1110001110110";
Trees_din <= "00000100000000000011110000001000";
wait for Clk_period;
Addr <= "1110001110111";
Trees_din <= "00000101000000000001100000000100";
wait for Clk_period;
Addr <= "1110001111000";
Trees_din <= "00000000001001010111001000010001";
wait for Clk_period;
Addr <= "1110001111001";
Trees_din <= "00000000001011110111001000010001";
wait for Clk_period;
Addr <= "1110001111010";
Trees_din <= "00000000000000000000011000000100";
wait for Clk_period;
Addr <= "1110001111011";
Trees_din <= "00000000000110110111001000010001";
wait for Clk_period;
Addr <= "1110001111100";
Trees_din <= "00000000000101000111001000010001";
wait for Clk_period;
Addr <= "1110001111101";
Trees_din <= "00000001000000000001101100001000";
wait for Clk_period;
Addr <= "1110001111110";
Trees_din <= "00000000000000000000101100000100";
wait for Clk_period;
Addr <= "1110001111111";
Trees_din <= "00000000010100100111001000010001";
wait for Clk_period;
Addr <= "1110010000000";
Trees_din <= "00000000000100110111001000010001";
wait for Clk_period;
Addr <= "1110010000001";
Trees_din <= "00000010000000000101110100000100";
wait for Clk_period;
Addr <= "1110010000010";
Trees_din <= "00000000010001100111001000010001";
wait for Clk_period;
Addr <= "1110010000011";
Trees_din <= "00000000000001110111001000010001";
wait for Clk_period;



----------tree 57-------------------

Addr <= "1110010000100";
Trees_din <= "00000101000000000010110010000000";
wait for Clk_period;
Addr <= "1110010000101";
Trees_din <= "00000010000000000000110101000000";
wait for Clk_period;
Addr <= "1110010000110";
Trees_din <= "00000001000000000001011000100000";
wait for Clk_period;
Addr <= "1110010000111";
Trees_din <= "00000001000000000001111100010000";
wait for Clk_period;
Addr <= "1110010001000";
Trees_din <= "00000110000000000010010100001000";
wait for Clk_period;
Addr <= "1110010001001";
Trees_din <= "00000101000000000011110000000100";
wait for Clk_period;
Addr <= "1110010001010";
Trees_din <= "00000000010100100111010000001101";
wait for Clk_period;
Addr <= "1110010001011";
Trees_din <= "00000000010000110111010000001101";
wait for Clk_period;
Addr <= "1110010001100";
Trees_din <= "00000010000000000001111000000100";
wait for Clk_period;
Addr <= "1110010001101";
Trees_din <= "00000000001100110111010000001101";
wait for Clk_period;
Addr <= "1110010001110";
Trees_din <= "00000000010000110111010000001101";
wait for Clk_period;
Addr <= "1110010001111";
Trees_din <= "00000010000000000101111100001000";
wait for Clk_period;
Addr <= "1110010010000";
Trees_din <= "00000011000000000010010000000100";
wait for Clk_period;
Addr <= "1110010010001";
Trees_din <= "00000000000101110111010000001101";
wait for Clk_period;
Addr <= "1110010010010";
Trees_din <= "00000000010100100111010000001101";
wait for Clk_period;
Addr <= "1110010010011";
Trees_din <= "00000001000000000001111000000100";
wait for Clk_period;
Addr <= "1110010010100";
Trees_din <= "00000000000100010111010000001101";
wait for Clk_period;
Addr <= "1110010010101";
Trees_din <= "00000000001100100111010000001101";
wait for Clk_period;
Addr <= "1110010010110";
Trees_din <= "00000111000000000011100000010000";
wait for Clk_period;
Addr <= "1110010010111";
Trees_din <= "00000000000000000001010100001000";
wait for Clk_period;
Addr <= "1110010011000";
Trees_din <= "00000111000000000000101000000100";
wait for Clk_period;
Addr <= "1110010011001";
Trees_din <= "00000000010110110111010000001101";
wait for Clk_period;
Addr <= "1110010011010";
Trees_din <= "00000000010111010111010000001101";
wait for Clk_period;
Addr <= "1110010011011";
Trees_din <= "00000110000000000100101000000100";
wait for Clk_period;
Addr <= "1110010011100";
Trees_din <= "00000000010101000111010000001101";
wait for Clk_period;
Addr <= "1110010011101";
Trees_din <= "00000000000000110111010000001101";
wait for Clk_period;
Addr <= "1110010011110";
Trees_din <= "00000000000000000100010100001000";
wait for Clk_period;
Addr <= "1110010011111";
Trees_din <= "00000010000000000101111100000100";
wait for Clk_period;
Addr <= "1110010100000";
Trees_din <= "00000000010010110111010000001101";
wait for Clk_period;
Addr <= "1110010100001";
Trees_din <= "00000000010100000111010000001101";
wait for Clk_period;
Addr <= "1110010100010";
Trees_din <= "00000001000000000010111000000100";
wait for Clk_period;
Addr <= "1110010100011";
Trees_din <= "00000000001100100111010000001101";
wait for Clk_period;
Addr <= "1110010100100";
Trees_din <= "00000000000101110111010000001101";
wait for Clk_period;
Addr <= "1110010100101";
Trees_din <= "00000011000000000000001000100000";
wait for Clk_period;
Addr <= "1110010100110";
Trees_din <= "00000100000000000000111100010000";
wait for Clk_period;
Addr <= "1110010100111";
Trees_din <= "00000010000000000011010100001000";
wait for Clk_period;
Addr <= "1110010101000";
Trees_din <= "00000000000000000010011000000100";
wait for Clk_period;
Addr <= "1110010101001";
Trees_din <= "00000000010011100111010000001101";
wait for Clk_period;
Addr <= "1110010101010";
Trees_din <= "00000000010011010111010000001101";
wait for Clk_period;
Addr <= "1110010101011";
Trees_din <= "00000010000000000101001100000100";
wait for Clk_period;
Addr <= "1110010101100";
Trees_din <= "00000000010101010111010000001101";
wait for Clk_period;
Addr <= "1110010101101";
Trees_din <= "00000000001010110111010000001101";
wait for Clk_period;
Addr <= "1110010101110";
Trees_din <= "00000110000000000110000100001000";
wait for Clk_period;
Addr <= "1110010101111";
Trees_din <= "00000010000000000100011100000100";
wait for Clk_period;
Addr <= "1110010110000";
Trees_din <= "00000000001011000111010000001101";
wait for Clk_period;
Addr <= "1110010110001";
Trees_din <= "00000000010011010111010000001101";
wait for Clk_period;
Addr <= "1110010110010";
Trees_din <= "00000001000000000100001100000100";
wait for Clk_period;
Addr <= "1110010110011";
Trees_din <= "00000000001111110111010000001101";
wait for Clk_period;
Addr <= "1110010110100";
Trees_din <= "00000000001000100111010000001101";
wait for Clk_period;
Addr <= "1110010110101";
Trees_din <= "00000000000000000100110000010000";
wait for Clk_period;
Addr <= "1110010110110";
Trees_din <= "00000000000000000001011100001000";
wait for Clk_period;
Addr <= "1110010110111";
Trees_din <= "00000010000000000010110000000100";
wait for Clk_period;
Addr <= "1110010111000";
Trees_din <= "00000000010101000111010000001101";
wait for Clk_period;
Addr <= "1110010111001";
Trees_din <= "00000000001001010111010000001101";
wait for Clk_period;
Addr <= "1110010111010";
Trees_din <= "00000011000000000011100100000100";
wait for Clk_period;
Addr <= "1110010111011";
Trees_din <= "00000000000111110111010000001101";
wait for Clk_period;
Addr <= "1110010111100";
Trees_din <= "00000000000000100111010000001101";
wait for Clk_period;
Addr <= "1110010111101";
Trees_din <= "00000100000000000011001100001000";
wait for Clk_period;
Addr <= "1110010111110";
Trees_din <= "00000001000000000001001000000100";
wait for Clk_period;
Addr <= "1110010111111";
Trees_din <= "00000000001110100111010000001101";
wait for Clk_period;
Addr <= "1110011000000";
Trees_din <= "00000000010100110111010000001101";
wait for Clk_period;
Addr <= "1110011000001";
Trees_din <= "00000001000000000000011000000100";
wait for Clk_period;
Addr <= "1110011000010";
Trees_din <= "00000000000000010111010000001101";
wait for Clk_period;
Addr <= "1110011000011";
Trees_din <= "00000000001101000111010000001101";
wait for Clk_period;
Addr <= "1110011000100";
Trees_din <= "00000100000000000100000101000000";
wait for Clk_period;
Addr <= "1110011000101";
Trees_din <= "00000110000000000011110100100000";
wait for Clk_period;
Addr <= "1110011000110";
Trees_din <= "00000110000000000100100100010000";
wait for Clk_period;
Addr <= "1110011000111";
Trees_din <= "00000011000000000100101000001000";
wait for Clk_period;
Addr <= "1110011001000";
Trees_din <= "00000101000000000000111000000100";
wait for Clk_period;
Addr <= "1110011001001";
Trees_din <= "00000000010110010111010000001101";
wait for Clk_period;
Addr <= "1110011001010";
Trees_din <= "00000000001110010111010000001101";
wait for Clk_period;
Addr <= "1110011001011";
Trees_din <= "00000000000000000010110000000100";
wait for Clk_period;
Addr <= "1110011001100";
Trees_din <= "00000000000010100111010000001101";
wait for Clk_period;
Addr <= "1110011001101";
Trees_din <= "00000000010001000111010000001101";
wait for Clk_period;
Addr <= "1110011001110";
Trees_din <= "00000000000000000010010000001000";
wait for Clk_period;
Addr <= "1110011001111";
Trees_din <= "00000100000000000101011100000100";
wait for Clk_period;
Addr <= "1110011010000";
Trees_din <= "00000000010010110111010000001101";
wait for Clk_period;
Addr <= "1110011010001";
Trees_din <= "00000000001111110111010000001101";
wait for Clk_period;
Addr <= "1110011010010";
Trees_din <= "00000100000000000101001100000100";
wait for Clk_period;
Addr <= "1110011010011";
Trees_din <= "00000000000111110111010000001101";
wait for Clk_period;
Addr <= "1110011010100";
Trees_din <= "00000000011000010111010000001101";
wait for Clk_period;
Addr <= "1110011010101";
Trees_din <= "00000101000000000101101000010000";
wait for Clk_period;
Addr <= "1110011010110";
Trees_din <= "00000000000000000000000100001000";
wait for Clk_period;
Addr <= "1110011010111";
Trees_din <= "00000001000000000001111100000100";
wait for Clk_period;
Addr <= "1110011011000";
Trees_din <= "00000000000000000111010000001101";
wait for Clk_period;
Addr <= "1110011011001";
Trees_din <= "00000000001101000111010000001101";
wait for Clk_period;
Addr <= "1110011011010";
Trees_din <= "00000100000000000010001000000100";
wait for Clk_period;
Addr <= "1110011011011";
Trees_din <= "00000000001010100111010000001101";
wait for Clk_period;
Addr <= "1110011011100";
Trees_din <= "00000000000111010111010000001101";
wait for Clk_period;
Addr <= "1110011011101";
Trees_din <= "00000100000000000101100100001000";
wait for Clk_period;
Addr <= "1110011011110";
Trees_din <= "00000111000000000011101100000100";
wait for Clk_period;
Addr <= "1110011011111";
Trees_din <= "00000000011000100111010000001101";
wait for Clk_period;
Addr <= "1110011100000";
Trees_din <= "00000000010010100111010000001101";
wait for Clk_period;
Addr <= "1110011100001";
Trees_din <= "00000010000000000100010100000100";
wait for Clk_period;
Addr <= "1110011100010";
Trees_din <= "00000000001110000111010000001101";
wait for Clk_period;
Addr <= "1110011100011";
Trees_din <= "00000000000110110111010000001101";
wait for Clk_period;
Addr <= "1110011100100";
Trees_din <= "00000100000000000110000100100000";
wait for Clk_period;
Addr <= "1110011100101";
Trees_din <= "00000100000000000100111000010000";
wait for Clk_period;
Addr <= "1110011100110";
Trees_din <= "00000010000000000101000000001000";
wait for Clk_period;
Addr <= "1110011100111";
Trees_din <= "00000101000000000011110100000100";
wait for Clk_period;
Addr <= "1110011101000";
Trees_din <= "00000000010111000111010000001101";
wait for Clk_period;
Addr <= "1110011101001";
Trees_din <= "00000000001011000111010000001101";
wait for Clk_period;
Addr <= "1110011101010";
Trees_din <= "00000111000000000011100100000100";
wait for Clk_period;
Addr <= "1110011101011";
Trees_din <= "00000000001000000111010000001101";
wait for Clk_period;
Addr <= "1110011101100";
Trees_din <= "00000000001111000111010000001101";
wait for Clk_period;
Addr <= "1110011101101";
Trees_din <= "00000000000000000011000100001000";
wait for Clk_period;
Addr <= "1110011101110";
Trees_din <= "00000011000000000101111000000100";
wait for Clk_period;
Addr <= "1110011101111";
Trees_din <= "00000000001010110111010000001101";
wait for Clk_period;
Addr <= "1110011110000";
Trees_din <= "00000000001000100111010000001101";
wait for Clk_period;
Addr <= "1110011110001";
Trees_din <= "00000110000000000000101100000100";
wait for Clk_period;
Addr <= "1110011110010";
Trees_din <= "00000000001110010111010000001101";
wait for Clk_period;
Addr <= "1110011110011";
Trees_din <= "00000000010110000111010000001101";
wait for Clk_period;
Addr <= "1110011110100";
Trees_din <= "00000101000000000100010000010000";
wait for Clk_period;
Addr <= "1110011110101";
Trees_din <= "00000100000000000011011000001000";
wait for Clk_period;
Addr <= "1110011110110";
Trees_din <= "00000101000000000011100100000100";
wait for Clk_period;
Addr <= "1110011110111";
Trees_din <= "00000000000111110111010000001101";
wait for Clk_period;
Addr <= "1110011111000";
Trees_din <= "00000000010101000111010000001101";
wait for Clk_period;
Addr <= "1110011111001";
Trees_din <= "00000001000000000101110000000100";
wait for Clk_period;
Addr <= "1110011111010";
Trees_din <= "00000000001101100111010000001101";
wait for Clk_period;
Addr <= "1110011111011";
Trees_din <= "00000000010011110111010000001101";
wait for Clk_period;
Addr <= "1110011111100";
Trees_din <= "00000100000000000001011100001000";
wait for Clk_period;
Addr <= "1110011111101";
Trees_din <= "00000001000000000100011000000100";
wait for Clk_period;
Addr <= "1110011111110";
Trees_din <= "00000000001000100111010000001101";
wait for Clk_period;
Addr <= "1110011111111";
Trees_din <= "00000000001100100111010000001101";
wait for Clk_period;
Addr <= "1110100000000";
Trees_din <= "00000011000000000010111100000100";
wait for Clk_period;
Addr <= "1110100000001";
Trees_din <= "00000000010000100111010000001101";
wait for Clk_period;
Addr <= "1110100000010";
Trees_din <= "00000000001101010111010000001101";
wait for Clk_period;



----------tree 58-------------------

Addr <= "1110100000011";
Trees_din <= "00000000000000000000111110000000";
wait for Clk_period;
Addr <= "1110100000100";
Trees_din <= "00000000000000000011000101000000";
wait for Clk_period;
Addr <= "1110100000101";
Trees_din <= "00000110000000000000010100100000";
wait for Clk_period;
Addr <= "1110100000110";
Trees_din <= "00000111000000000000000100010000";
wait for Clk_period;
Addr <= "1110100000111";
Trees_din <= "00000111000000000000011000001000";
wait for Clk_period;
Addr <= "1110100001000";
Trees_din <= "00000100000000000010010000000100";
wait for Clk_period;
Addr <= "1110100001001";
Trees_din <= "00000000001011000111011000001001";
wait for Clk_period;
Addr <= "1110100001010";
Trees_din <= "00000000001101000111011000001001";
wait for Clk_period;
Addr <= "1110100001011";
Trees_din <= "00000011000000000101101100000100";
wait for Clk_period;
Addr <= "1110100001100";
Trees_din <= "00000000000100100111011000001001";
wait for Clk_period;
Addr <= "1110100001101";
Trees_din <= "00000000010100100111011000001001";
wait for Clk_period;
Addr <= "1110100001110";
Trees_din <= "00000010000000000010101100001000";
wait for Clk_period;
Addr <= "1110100001111";
Trees_din <= "00000011000000000010010100000100";
wait for Clk_period;
Addr <= "1110100010000";
Trees_din <= "00000000001100000111011000001001";
wait for Clk_period;
Addr <= "1110100010001";
Trees_din <= "00000000000110110111011000001001";
wait for Clk_period;
Addr <= "1110100010010";
Trees_din <= "00000111000000000010011000000100";
wait for Clk_period;
Addr <= "1110100010011";
Trees_din <= "00000000011000010111011000001001";
wait for Clk_period;
Addr <= "1110100010100";
Trees_din <= "00000000001001110111011000001001";
wait for Clk_period;
Addr <= "1110100010101";
Trees_din <= "00000000000000000101111000010000";
wait for Clk_period;
Addr <= "1110100010110";
Trees_din <= "00000111000000000000100000001000";
wait for Clk_period;
Addr <= "1110100010111";
Trees_din <= "00000110000000000100011100000100";
wait for Clk_period;
Addr <= "1110100011000";
Trees_din <= "00000000010110000111011000001001";
wait for Clk_period;
Addr <= "1110100011001";
Trees_din <= "00000000010011110111011000001001";
wait for Clk_period;
Addr <= "1110100011010";
Trees_din <= "00000011000000000011000100000100";
wait for Clk_period;
Addr <= "1110100011011";
Trees_din <= "00000000001011010111011000001001";
wait for Clk_period;
Addr <= "1110100011100";
Trees_din <= "00000000000111010111011000001001";
wait for Clk_period;
Addr <= "1110100011101";
Trees_din <= "00000001000000000101000100001000";
wait for Clk_period;
Addr <= "1110100011110";
Trees_din <= "00000011000000000010010100000100";
wait for Clk_period;
Addr <= "1110100011111";
Trees_din <= "00000000010110010111011000001001";
wait for Clk_period;
Addr <= "1110100100000";
Trees_din <= "00000000001011010111011000001001";
wait for Clk_period;
Addr <= "1110100100001";
Trees_din <= "00000000000000000011000000000100";
wait for Clk_period;
Addr <= "1110100100010";
Trees_din <= "00000000000110000111011000001001";
wait for Clk_period;
Addr <= "1110100100011";
Trees_din <= "00000000001010100111011000001001";
wait for Clk_period;
Addr <= "1110100100100";
Trees_din <= "00000001000000000000100100100000";
wait for Clk_period;
Addr <= "1110100100101";
Trees_din <= "00000000000000000000111000010000";
wait for Clk_period;
Addr <= "1110100100110";
Trees_din <= "00000011000000000101101100001000";
wait for Clk_period;
Addr <= "1110100100111";
Trees_din <= "00000110000000000011111000000100";
wait for Clk_period;
Addr <= "1110100101000";
Trees_din <= "00000000000001000111011000001001";
wait for Clk_period;
Addr <= "1110100101001";
Trees_din <= "00000000001111000111011000001001";
wait for Clk_period;
Addr <= "1110100101010";
Trees_din <= "00000011000000000100011100000100";
wait for Clk_period;
Addr <= "1110100101011";
Trees_din <= "00000000011000010111011000001001";
wait for Clk_period;
Addr <= "1110100101100";
Trees_din <= "00000000011000100111011000001001";
wait for Clk_period;
Addr <= "1110100101101";
Trees_din <= "00000011000000000010111000001000";
wait for Clk_period;
Addr <= "1110100101110";
Trees_din <= "00000101000000000001001000000100";
wait for Clk_period;
Addr <= "1110100101111";
Trees_din <= "00000000000110010111011000001001";
wait for Clk_period;
Addr <= "1110100110000";
Trees_din <= "00000000001000110111011000001001";
wait for Clk_period;
Addr <= "1110100110001";
Trees_din <= "00000110000000000000100000000100";
wait for Clk_period;
Addr <= "1110100110010";
Trees_din <= "00000000001101000111011000001001";
wait for Clk_period;
Addr <= "1110100110011";
Trees_din <= "00000000001110010111011000001001";
wait for Clk_period;
Addr <= "1110100110100";
Trees_din <= "00000000000000000011001000010000";
wait for Clk_period;
Addr <= "1110100110101";
Trees_din <= "00000100000000000100110100001000";
wait for Clk_period;
Addr <= "1110100110110";
Trees_din <= "00000010000000000001111000000100";
wait for Clk_period;
Addr <= "1110100110111";
Trees_din <= "00000000000101010111011000001001";
wait for Clk_period;
Addr <= "1110100111000";
Trees_din <= "00000000010100000111011000001001";
wait for Clk_period;
Addr <= "1110100111001";
Trees_din <= "00000101000000000000011000000100";
wait for Clk_period;
Addr <= "1110100111010";
Trees_din <= "00000000000111110111011000001001";
wait for Clk_period;
Addr <= "1110100111011";
Trees_din <= "00000000001010000111011000001001";
wait for Clk_period;
Addr <= "1110100111100";
Trees_din <= "00000011000000000010110000001000";
wait for Clk_period;
Addr <= "1110100111101";
Trees_din <= "00000010000000000110001100000100";
wait for Clk_period;
Addr <= "1110100111110";
Trees_din <= "00000000000010110111011000001001";
wait for Clk_period;
Addr <= "1110100111111";
Trees_din <= "00000000001000110111011000001001";
wait for Clk_period;
Addr <= "1110101000000";
Trees_din <= "00000001000000000100000000000100";
wait for Clk_period;
Addr <= "1110101000001";
Trees_din <= "00000000010011110111011000001001";
wait for Clk_period;
Addr <= "1110101000010";
Trees_din <= "00000000001001000111011000001001";
wait for Clk_period;
Addr <= "1110101000011";
Trees_din <= "00000010000000000011111101000000";
wait for Clk_period;
Addr <= "1110101000100";
Trees_din <= "00000101000000000011101000100000";
wait for Clk_period;
Addr <= "1110101000101";
Trees_din <= "00000000000000000001111000010000";
wait for Clk_period;
Addr <= "1110101000110";
Trees_din <= "00000100000000000101000000001000";
wait for Clk_period;
Addr <= "1110101000111";
Trees_din <= "00000111000000000000001100000100";
wait for Clk_period;
Addr <= "1110101001000";
Trees_din <= "00000000011001000111011000001001";
wait for Clk_period;
Addr <= "1110101001001";
Trees_din <= "00000000001010110111011000001001";
wait for Clk_period;
Addr <= "1110101001010";
Trees_din <= "00000001000000000001110100000100";
wait for Clk_period;
Addr <= "1110101001011";
Trees_din <= "00000000010101000111011000001001";
wait for Clk_period;
Addr <= "1110101001100";
Trees_din <= "00000000010111000111011000001001";
wait for Clk_period;
Addr <= "1110101001101";
Trees_din <= "00000100000000000010111000001000";
wait for Clk_period;
Addr <= "1110101001110";
Trees_din <= "00000011000000000100011000000100";
wait for Clk_period;
Addr <= "1110101001111";
Trees_din <= "00000000010001010111011000001001";
wait for Clk_period;
Addr <= "1110101010000";
Trees_din <= "00000000000110000111011000001001";
wait for Clk_period;
Addr <= "1110101010001";
Trees_din <= "00000011000000000101011000000100";
wait for Clk_period;
Addr <= "1110101010010";
Trees_din <= "00000000010101000111011000001001";
wait for Clk_period;
Addr <= "1110101010011";
Trees_din <= "00000000001110100111011000001001";
wait for Clk_period;
Addr <= "1110101010100";
Trees_din <= "00000011000000000100110100010000";
wait for Clk_period;
Addr <= "1110101010101";
Trees_din <= "00000100000000000001111100001000";
wait for Clk_period;
Addr <= "1110101010110";
Trees_din <= "00000100000000000101000000000100";
wait for Clk_period;
Addr <= "1110101010111";
Trees_din <= "00000000010100110111011000001001";
wait for Clk_period;
Addr <= "1110101011000";
Trees_din <= "00000000001011110111011000001001";
wait for Clk_period;
Addr <= "1110101011001";
Trees_din <= "00000011000000000001000000000100";
wait for Clk_period;
Addr <= "1110101011010";
Trees_din <= "00000000010001100111011000001001";
wait for Clk_period;
Addr <= "1110101011011";
Trees_din <= "00000000001010010111011000001001";
wait for Clk_period;
Addr <= "1110101011100";
Trees_din <= "00000011000000000001010100001000";
wait for Clk_period;
Addr <= "1110101011101";
Trees_din <= "00000001000000000010001000000100";
wait for Clk_period;
Addr <= "1110101011110";
Trees_din <= "00000000010001000111011000001001";
wait for Clk_period;
Addr <= "1110101011111";
Trees_din <= "00000000001000100111011000001001";
wait for Clk_period;
Addr <= "1110101100000";
Trees_din <= "00000001000000000010011100000100";
wait for Clk_period;
Addr <= "1110101100001";
Trees_din <= "00000000000011100111011000001001";
wait for Clk_period;
Addr <= "1110101100010";
Trees_din <= "00000000000001110111011000001001";
wait for Clk_period;
Addr <= "1110101100011";
Trees_din <= "00000000000000000100001000100000";
wait for Clk_period;
Addr <= "1110101100100";
Trees_din <= "00000011000000000110001100010000";
wait for Clk_period;
Addr <= "1110101100101";
Trees_din <= "00000001000000000011000100001000";
wait for Clk_period;
Addr <= "1110101100110";
Trees_din <= "00000110000000000000000100000100";
wait for Clk_period;
Addr <= "1110101100111";
Trees_din <= "00000000001001010111011000001001";
wait for Clk_period;
Addr <= "1110101101000";
Trees_din <= "00000000010011010111011000001001";
wait for Clk_period;
Addr <= "1110101101001";
Trees_din <= "00000101000000000001000000000100";
wait for Clk_period;
Addr <= "1110101101010";
Trees_din <= "00000000001100110111011000001001";
wait for Clk_period;
Addr <= "1110101101011";
Trees_din <= "00000000010011100111011000001001";
wait for Clk_period;
Addr <= "1110101101100";
Trees_din <= "00000010000000000011001100001000";
wait for Clk_period;
Addr <= "1110101101101";
Trees_din <= "00000111000000000100011000000100";
wait for Clk_period;
Addr <= "1110101101110";
Trees_din <= "00000000000100000111011000001001";
wait for Clk_period;
Addr <= "1110101101111";
Trees_din <= "00000000001110100111011000001001";
wait for Clk_period;
Addr <= "1110101110000";
Trees_din <= "00000101000000000001100000000100";
wait for Clk_period;
Addr <= "1110101110001";
Trees_din <= "00000000001110100111011000001001";
wait for Clk_period;
Addr <= "1110101110010";
Trees_din <= "00000000011000010111011000001001";
wait for Clk_period;
Addr <= "1110101110011";
Trees_din <= "00000000000000000011101100010000";
wait for Clk_period;
Addr <= "1110101110100";
Trees_din <= "00000001000000000000110000001000";
wait for Clk_period;
Addr <= "1110101110101";
Trees_din <= "00000010000000000110010000000100";
wait for Clk_period;
Addr <= "1110101110110";
Trees_din <= "00000000001000000111011000001001";
wait for Clk_period;
Addr <= "1110101110111";
Trees_din <= "00000000010100010111011000001001";
wait for Clk_period;
Addr <= "1110101111000";
Trees_din <= "00000101000000000011101100000100";
wait for Clk_period;
Addr <= "1110101111001";
Trees_din <= "00000000001100010111011000001001";
wait for Clk_period;
Addr <= "1110101111010";
Trees_din <= "00000000010001000111011000001001";
wait for Clk_period;
Addr <= "1110101111011";
Trees_din <= "00000001000000000110001100001000";
wait for Clk_period;
Addr <= "1110101111100";
Trees_din <= "00000101000000000110000000000100";
wait for Clk_period;
Addr <= "1110101111101";
Trees_din <= "00000000000100010111011000001001";
wait for Clk_period;
Addr <= "1110101111110";
Trees_din <= "00000000001100110111011000001001";
wait for Clk_period;
Addr <= "1110101111111";
Trees_din <= "00000101000000000000000000000100";
wait for Clk_period;
Addr <= "1110110000000";
Trees_din <= "00000000000010100111011000001001";
wait for Clk_period;
Addr <= "1110110000001";
Trees_din <= "00000000010010000111011000001001";
wait for Clk_period;



----------tree 59-------------------

Addr <= "1110110000010";
Trees_din <= "00000110000000000001111110000000";
wait for Clk_period;
Addr <= "1110110000011";
Trees_din <= "00000111000000000010010001000000";
wait for Clk_period;
Addr <= "1110110000100";
Trees_din <= "00000101000000000101100100100000";
wait for Clk_period;
Addr <= "1110110000101";
Trees_din <= "00000111000000000010110100010000";
wait for Clk_period;
Addr <= "1110110000110";
Trees_din <= "00000100000000000101100000001000";
wait for Clk_period;
Addr <= "1110110000111";
Trees_din <= "00000010000000000001100000000100";
wait for Clk_period;
Addr <= "1110110001000";
Trees_din <= "00000000010010110000000000000011";
wait for Clk_period;
Addr <= "1110110001001";
Trees_din <= "00000000000110110000000000000011";
wait for Clk_period;
Addr <= "1110110001010";
Trees_din <= "00000000000000000011100000000100";
wait for Clk_period;
Addr <= "1110110001011";
Trees_din <= "00000000010110110000000000000011";
wait for Clk_period;
Addr <= "1110110001100";
Trees_din <= "00000000010110110000000000000011";
wait for Clk_period;
Addr <= "1110110001101";
Trees_din <= "00000001000000000110000000001000";
wait for Clk_period;
Addr <= "1110110001110";
Trees_din <= "00000001000000000100000000000100";
wait for Clk_period;
Addr <= "1110110001111";
Trees_din <= "00000000000101000000000000000011";
wait for Clk_period;
Addr <= "1110110010000";
Trees_din <= "00000000001111010000000000000011";
wait for Clk_period;
Addr <= "1110110010001";
Trees_din <= "00000100000000000001111100000100";
wait for Clk_period;
Addr <= "1110110010010";
Trees_din <= "00000000001110010000000000000011";
wait for Clk_period;
Addr <= "1110110010011";
Trees_din <= "00000000010101010000000000000011";
wait for Clk_period;
Addr <= "1110110010100";
Trees_din <= "00000011000000000100010000010000";
wait for Clk_period;
Addr <= "1110110010101";
Trees_din <= "00000011000000000100110100001000";
wait for Clk_period;
Addr <= "1110110010110";
Trees_din <= "00000101000000000101001100000100";
wait for Clk_period;
Addr <= "1110110010111";
Trees_din <= "00000000000001100000000000000011";
wait for Clk_period;
Addr <= "1110110011000";
Trees_din <= "00000000000011000000000000000011";
wait for Clk_period;
Addr <= "1110110011001";
Trees_din <= "00000010000000000010000100000100";
wait for Clk_period;
Addr <= "1110110011010";
Trees_din <= "00000000001010010000000000000011";
wait for Clk_period;
Addr <= "1110110011011";
Trees_din <= "00000000001100010000000000000011";
wait for Clk_period;
Addr <= "1110110011100";
Trees_din <= "00000111000000000100111100001000";
wait for Clk_period;
Addr <= "1110110011101";
Trees_din <= "00000000000000000100111100000100";
wait for Clk_period;
Addr <= "1110110011110";
Trees_din <= "00000000000001110000000000000011";
wait for Clk_period;
Addr <= "1110110011111";
Trees_din <= "00000000001101000000000000000011";
wait for Clk_period;
Addr <= "1110110100000";
Trees_din <= "00000011000000000001011100000100";
wait for Clk_period;
Addr <= "1110110100001";
Trees_din <= "00000000001000110000000000000011";
wait for Clk_period;
Addr <= "1110110100010";
Trees_din <= "00000000001101010000000000000011";
wait for Clk_period;
Addr <= "1110110100011";
Trees_din <= "00000101000000000101001100100000";
wait for Clk_period;
Addr <= "1110110100100";
Trees_din <= "00000111000000000010001100010000";
wait for Clk_period;
Addr <= "1110110100101";
Trees_din <= "00000111000000000101001100001000";
wait for Clk_period;
Addr <= "1110110100110";
Trees_din <= "00000000000000000011101100000100";
wait for Clk_period;
Addr <= "1110110100111";
Trees_din <= "00000000001101000000000000000011";
wait for Clk_period;
Addr <= "1110110101000";
Trees_din <= "00000000010110100000000000000011";
wait for Clk_period;
Addr <= "1110110101001";
Trees_din <= "00000101000000000011110000000100";
wait for Clk_period;
Addr <= "1110110101010";
Trees_din <= "00000000000010010000000000000011";
wait for Clk_period;
Addr <= "1110110101011";
Trees_din <= "00000000010110010000000000000011";
wait for Clk_period;
Addr <= "1110110101100";
Trees_din <= "00000100000000000101010100001000";
wait for Clk_period;
Addr <= "1110110101101";
Trees_din <= "00000100000000000010001000000100";
wait for Clk_period;
Addr <= "1110110101110";
Trees_din <= "00000000011000000000000000000011";
wait for Clk_period;
Addr <= "1110110101111";
Trees_din <= "00000000001111000000000000000011";
wait for Clk_period;
Addr <= "1110110110000";
Trees_din <= "00000100000000000000000100000100";
wait for Clk_period;
Addr <= "1110110110001";
Trees_din <= "00000000001101100000000000000011";
wait for Clk_period;
Addr <= "1110110110010";
Trees_din <= "00000000010110000000000000000011";
wait for Clk_period;
Addr <= "1110110110011";
Trees_din <= "00000001000000000011110100010000";
wait for Clk_period;
Addr <= "1110110110100";
Trees_din <= "00000101000000000100111100001000";
wait for Clk_period;
Addr <= "1110110110101";
Trees_din <= "00000100000000000100111100000100";
wait for Clk_period;
Addr <= "1110110110110";
Trees_din <= "00000000000101110000000000000011";
wait for Clk_period;
Addr <= "1110110110111";
Trees_din <= "00000000000101010000000000000011";
wait for Clk_period;
Addr <= "1110110111000";
Trees_din <= "00000110000000000101100000000100";
wait for Clk_period;
Addr <= "1110110111001";
Trees_din <= "00000000000001110000000000000011";
wait for Clk_period;
Addr <= "1110110111010";
Trees_din <= "00000000011000100000000000000011";
wait for Clk_period;
Addr <= "1110110111011";
Trees_din <= "00000000000000000100111100001000";
wait for Clk_period;
Addr <= "1110110111100";
Trees_din <= "00000001000000000001001100000100";
wait for Clk_period;
Addr <= "1110110111101";
Trees_din <= "00000000001011010000000000000011";
wait for Clk_period;
Addr <= "1110110111110";
Trees_din <= "00000000001101010000000000000011";
wait for Clk_period;
Addr <= "1110110111111";
Trees_din <= "00000010000000000100111000000100";
wait for Clk_period;
Addr <= "1110111000000";
Trees_din <= "00000000000011010000000000000011";
wait for Clk_period;
Addr <= "1110111000001";
Trees_din <= "00000000010010000000000000000011";
wait for Clk_period;
Addr <= "1110111000010";
Trees_din <= "00000000000000000101000101000000";
wait for Clk_period;
Addr <= "1110111000011";
Trees_din <= "00000011000000000101010000100000";
wait for Clk_period;
Addr <= "1110111000100";
Trees_din <= "00000000000000000010010000010000";
wait for Clk_period;
Addr <= "1110111000101";
Trees_din <= "00000111000000000010101000001000";
wait for Clk_period;
Addr <= "1110111000110";
Trees_din <= "00000110000000000000001000000100";
wait for Clk_period;
Addr <= "1110111000111";
Trees_din <= "00000000001101010000000000000011";
wait for Clk_period;
Addr <= "1110111001000";
Trees_din <= "00000000010001100000000000000011";
wait for Clk_period;
Addr <= "1110111001001";
Trees_din <= "00000101000000000101101000000100";
wait for Clk_period;
Addr <= "1110111001010";
Trees_din <= "00000000001010110000000000000011";
wait for Clk_period;
Addr <= "1110111001011";
Trees_din <= "00000000001100100000000000000011";
wait for Clk_period;
Addr <= "1110111001100";
Trees_din <= "00000110000000000010001100001000";
wait for Clk_period;
Addr <= "1110111001101";
Trees_din <= "00000111000000000101100000000100";
wait for Clk_period;
Addr <= "1110111001110";
Trees_din <= "00000000001110100000000000000011";
wait for Clk_period;
Addr <= "1110111001111";
Trees_din <= "00000000001110100000000000000011";
wait for Clk_period;
Addr <= "1110111010000";
Trees_din <= "00000011000000000001000000000100";
wait for Clk_period;
Addr <= "1110111010001";
Trees_din <= "00000000010001000000000000000011";
wait for Clk_period;
Addr <= "1110111010010";
Trees_din <= "00000000001001010000000000000011";
wait for Clk_period;
Addr <= "1110111010011";
Trees_din <= "00000011000000000011110000010000";
wait for Clk_period;
Addr <= "1110111010100";
Trees_din <= "00000010000000000010111100001000";
wait for Clk_period;
Addr <= "1110111010101";
Trees_din <= "00000011000000000110000000000100";
wait for Clk_period;
Addr <= "1110111010110";
Trees_din <= "00000000000100010000000000000011";
wait for Clk_period;
Addr <= "1110111010111";
Trees_din <= "00000000000001100000000000000011";
wait for Clk_period;
Addr <= "1110111011000";
Trees_din <= "00000110000000000011000100000100";
wait for Clk_period;
Addr <= "1110111011001";
Trees_din <= "00000000011001000000000000000011";
wait for Clk_period;
Addr <= "1110111011010";
Trees_din <= "00000000001111110000000000000011";
wait for Clk_period;
Addr <= "1110111011011";
Trees_din <= "00000100000000000100110100001000";
wait for Clk_period;
Addr <= "1110111011100";
Trees_din <= "00000010000000000011100100000100";
wait for Clk_period;
Addr <= "1110111011101";
Trees_din <= "00000000000100010000000000000011";
wait for Clk_period;
Addr <= "1110111011110";
Trees_din <= "00000000000001000000000000000011";
wait for Clk_period;
Addr <= "1110111011111";
Trees_din <= "00000100000000000000000100000100";
wait for Clk_period;
Addr <= "1110111100000";
Trees_din <= "00000000001010100000000000000011";
wait for Clk_period;
Addr <= "1110111100001";
Trees_din <= "00000000010000100000000000000011";
wait for Clk_period;
Addr <= "1110111100010";
Trees_din <= "00000101000000000011010000100000";
wait for Clk_period;
Addr <= "1110111100011";
Trees_din <= "00000000000000000100010000010000";
wait for Clk_period;
Addr <= "1110111100100";
Trees_din <= "00000101000000000100101100001000";
wait for Clk_period;
Addr <= "1110111100101";
Trees_din <= "00000101000000000101110100000100";
wait for Clk_period;
Addr <= "1110111100110";
Trees_din <= "00000000001010010000000000000011";
wait for Clk_period;
Addr <= "1110111100111";
Trees_din <= "00000000000001010000000000000011";
wait for Clk_period;
Addr <= "1110111101000";
Trees_din <= "00000010000000000011000100000100";
wait for Clk_period;
Addr <= "1110111101001";
Trees_din <= "00000000001000110000000000000011";
wait for Clk_period;
Addr <= "1110111101010";
Trees_din <= "00000000001110110000000000000011";
wait for Clk_period;
Addr <= "1110111101011";
Trees_din <= "00000100000000000010111000001000";
wait for Clk_period;
Addr <= "1110111101100";
Trees_din <= "00000100000000000011111100000100";
wait for Clk_period;
Addr <= "1110111101101";
Trees_din <= "00000000001100000000000000000011";
wait for Clk_period;
Addr <= "1110111101110";
Trees_din <= "00000000010001110000000000000011";
wait for Clk_period;
Addr <= "1110111101111";
Trees_din <= "00000111000000000001110100000100";
wait for Clk_period;
Addr <= "1110111110000";
Trees_din <= "00000000010000010000000000000011";
wait for Clk_period;
Addr <= "1110111110001";
Trees_din <= "00000000001001100000000000000011";
wait for Clk_period;
Addr <= "1110111110010";
Trees_din <= "00000100000000000100100000010000";
wait for Clk_period;
Addr <= "1110111110011";
Trees_din <= "00000001000000000000110100001000";
wait for Clk_period;
Addr <= "1110111110100";
Trees_din <= "00000110000000000100010000000100";
wait for Clk_period;
Addr <= "1110111110101";
Trees_din <= "00000000001110110000000000000011";
wait for Clk_period;
Addr <= "1110111110110";
Trees_din <= "00000000001101100000000000000011";
wait for Clk_period;
Addr <= "1110111110111";
Trees_din <= "00000111000000000100000000000100";
wait for Clk_period;
Addr <= "1110111111000";
Trees_din <= "00000000000110110000000000000011";
wait for Clk_period;
Addr <= "1110111111001";
Trees_din <= "00000000010110010000000000000011";
wait for Clk_period;
Addr <= "1110111111010";
Trees_din <= "00000111000000000010001000001000";
wait for Clk_period;
Addr <= "1110111111011";
Trees_din <= "00000011000000000001001000000100";
wait for Clk_period;
Addr <= "1110111111100";
Trees_din <= "00000000000101010000000000000011";
wait for Clk_period;
Addr <= "1110111111101";
Trees_din <= "00000000000010000000000000000011";
wait for Clk_period;
Addr <= "1110111111110";
Trees_din <= "00000101000000000010011100000100";
wait for Clk_period;
Addr <= "1110111111111";
Trees_din <= "00000000010011010000000000000011";
wait for Clk_period;
Addr <= "1111000000000";
Trees_din <= "00000000001111010000000000000011";
wait for Clk_period;


-- LOAD TREES END
-----------------------------------------------------------------------

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period;

        -- class_label <= std_logic_vector(to_unsigned(0, class_label'length));

        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';

-- LOAD FEATURES START
-----------------------------------------------------------------------

        Features_din <= "0000000000110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';

        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;
        Features_din <= "0000000000110010";
        wait for Clk_period;

        Last_feature <= '1';
        pc_count     <= '1';
        Features_din <= "0000000000110010";
        wait for Clk_period;

-- LOAD FEATURES START
-----------------------------------------------------------------------

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';

        -- Wait until inference is complete
        v_TIME := now;
        wait until Finish = '1';
        v_TIME := now - V_TIME;
        report "Execution Time = " & time'image(v_TIME);

        wait for Clk_period * 1/2;

        if Dout = class_label then
            hc_count <= '1';
        end if;

        wait for Clk_period;
        hc_count <= '0';

        stop;
    end process;
end;
    